PK   '6X137=�	  2\     cirkitFile.json�\�o�8�W�W��I�����=�a�z�=$�AIT#�#�d�i���~���rl�tf6]Nbqf8~�8K�t��iEۙ�ӭ�	�@͂;ݕ�z|5�u�����N?�W�����`¢�h��J��E�ԅsL��"�Ҵ̲8ZD�������@SG����K�~J9�+#�Cm�2���ì�*1&ϔ���}zV����������3"X#J؁v . � .�D}E�'���"r�]$�4R���?$���C"���?$���C"�b^�;ݽ'w�&~�m��5Nu]B���0���T�+��^�D���Ɏ�8�*�(̳Ⱥ]�2�+��UV�V2.���^J�$�穤�+^@�R��J�<�����BN35f�`z�'���1{�<Mc����iw�+�e�~�ߢ�uz����� ��bEn��Jd+�YI�Hk���eD	����Jƃ�xue�b���_��/H3������b�A1�P02q0���ȃb�A1�yP�<(F��(�='2X�sۋ�ɏ�q.�=U1�r>��<������e+�'	+<���O�W��5�o̺�����ӭ ��bE�XQ,Vb+	����Jƃ:&��x�<� �����a�1�yP�L̃b�A1�yP�<(F#��ł��,��}�_�.(�D�n��r�N�_�j�D�n��y'�t+<���b��|�7��E]~��Y�Xwf�xX�{h��t��5�7c�7����]�ڷ�����y��1O�J��{��G9�Qz��'��y������t��bYF7�)¹�N�4ֹu������y�u�	"���[P���I�g���"��V��� ������ ����y�1���u��jû�mU���.�e��`L�G�� 껃Tt���G���#�1et	Q?%�gTtE��$�
Br��W�v��(�**�
K����D*o"�8�HD*��D�"�HD*��D�"QP�(^@�w�����]�}f�zc�_��]�}f�vn��7|K�~����ֻ���w�w���ݣ�=͂���t���r)��jt7��1�0��tPs����b�N�;�owc�N�(8Yp������� N���:t�4�i��@��NC81<��i����X�Y8���9��D�1��bs'�l���y���1���y�2�1k���U��	���8�X|���f��!��w__-un�nY���_���-�c�Mp܄�&<n�&q�$�M�q�^.ygt���s%�],�U�b�T�U&�!Ve�
�P'v�2�,8��b�.�ݭ��%KS�ם6y;"��o������҇�}0]_�������:�껺�l��{�ٵ΂/z�v����;�]7��$�������?����˕��+�}�Wu�4�k����L\�v 6��YW��ם�^r`,6�dS^b����خ�~�/�!$b��f�\f�����U�{Q�[Ȋ0��&Ҳ��0�\�+�J�t0م���_g�����)6��v�Y�v���7.�g��N��:ù�I����чx�"�-b��hԒ���o9���������u��� Jγ� �&�M0�MjA:�ɴ��֒�Z8��ZCxO�$8բ&u�N�����u8m�v@�u��_�u�} s1w��`��Ň�]{�ʢtc2��X�!JA�-Վ���Z�U�ŨCU�������*�TUD��2���/Á~�/D�iG`�$�x.�$�lK$3�2�4������4�Ms����R��b'�I7I��1�I�Z^��Z3%�yB�"x�f�1!�V�a6-�J� v�$1s�E�ؼd���,bc�TIX(C����*��J�\�$�#U����l��cs4��%�e�HOl4Es�{a�W��=���������u�˻�\;;�8�fv�����#�f�Y�T*��03X�"�2f�IY�
/�x��<�a��$�3 � �j��t�9���]7倞�}p-b*���MW�%0���X����K�^��ԟ%ٽ����컲�.�L��.��Й����6��qwp����M0�@v\��x��&��X���P7�ʡ��'���i�M�tS�~��隵�O>�ں�?��n�����&p����k�8�ڕ�zu�~��C��h9�� %�˥$�SR��r�ín'���i�ۧ���� �bd~�]�s ���Avv�.��gR�:��b!��N�=~5+>����%(�0��O�z��=i�$�d�I�R�	�E�S�RoEQ���.�/-E�j<;M�)?H�<���e�t�/�xՁ��E]@,��q�z͜o�Yg��s�8;���x��)ux��I����i�G�9�G~_!0ț4.��b 	���X��?N��~R�՝I IM h��� ��0#x�_�*�J%���$$~R���I Im ���r���]�������VÇ���]7k����כ����S��PK   '6X��(��8  �8  /   images/02932828-f6d4-4923-89fb-67d65ebd103a.png�8!ǉPNG

   IHDR   d   �   ���   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  8kIDATx���T����������tX�,�(HS�(c��5�ؒ�1&�3��&�F�1�?1Ѩ�1��i"(�.,�l�;���o�웶�]��|ٙw�}�s���<ߘ1cZ����&�x<��z���K\\�466JKK��=!!a��f���f�w||��{���!x�#��1��|>�< �\�r���>�v�q���͛eӦM2e����dܸq2l�0ٹs�����	��}�G�ĉ���J^y�)//��=�IIIr��'˜9s$%%E;�0ٺu��q��.�E�u�(<�]p�:,��g��:9##C$999�x�m۶Iqq���Yd��=z�̜9S���Z�߿����K����g��C9������'//���'�0s:T�-[�_�y��Jee�A<�~��f��ٳG.��2Y�~�����KlϧO�>2`� IKK3g�޽��555!�A��Ғ��w�O��Ө(P�6rݺu�t�Ґ���v��an�U�J�ٳ�lٲEv��%EEEf�u���Y����3�\\��� ���s�]�}�v�����3c�p�n�4i�2��Z���^�>r���J��/6���gAX��t�0ax�R�%J9�t�$(u���Pޚ�������_���:�\��B���w������a�\���ZxFvʆ��n6���q};Vw�%��W�^�JAAAȯ���S|���c�����#	z��!cǎ���z����iJ�=�!v�#F�xAW��M�� 7ʶ}�����o�'�|R=�P����
�%tvn1+Y������� �畕+W�"L�n�,�e���V�Q�������ؕ�;,11�E�[��r��p)�*�B	��-�N�����P�W���9~�m��N�ͼ�_�כ<���
-���?�8O���h��TU�.��w�q�lۺM�9��y�	RUY%wnO�
As��>عc��=�9����o��V`��+������J�,^ I	>y��G���e��r�7N�Q#�ˋ�?+�e%���$��		�fa(^���_���%�w����7r�5ט�7��>K�K6� H�6;D���}W^ye��gϖ;���S]q��΀Ҭʐ��������<�w���eM��*�q���Q�Ƀ�Յ���&3$>c��dű�;�H�lʢ��d᧋͹��\I���y���/iƙ��v�_�w�<5w����J��������7�IrS��Iz��́����n��{ｆ((ʶv*�W�=�c��y<�ET�3�^8X�A�W�ҴZ���:�h��47���5�����|��/���S��رn�(���o-N�#�:TD{P$��߷�rK���.�j�>S[[kvKT>j�js�bn��|<����5��Zb�(��s�D��Ǽb�]�yc�ӑyU����<+,�9cΫ�dT��?Z]ǹ�����;�4�n��V��+**233�#��i���|�8��$:�#���A %H��<T� ���Ȋ��KmE������"i�x%��@��;\�S�Ϯ�x�i�\�y� q���)��=���|�^�'i=�IF�A�OT6�����2���U��%ez��U��KL���C$C?]��MQ�G�EM��Ç������޽{�sss�a���)!��Y�Ǒ����=?p��G�e���u�1%T��Q5���]��SZ�S|2�~)���J�����LK���ee]��|��t7T
 �-�d�s7If�Qr�ٿG���mPB�{�ϲo���'�Jz��뽪*��I*<$���Ȁ����؅�����d�+wI��)2�?��l�����3Y������Œ���z�U5��a^�T��e��ߓ���"m[D��[�r�jY�R�}II�T�6��a]��t���O>	�!2����������<�4��q*�.S{dȼy��;J�/QJ������L헱��K��s�qSJFZ���`�������u�����oB�C]���RQ�.�L+�Aj���ŏ^#Ǐ��+�"#�$9)^�A�U�2��5r�_~*{t�#ξI�g�aW�W�H�����#��Z��m�+����3��"��d�jƏ�"%����ܵr��W�ލɘS�	��V����by���� /��1N�����0���s�ƍ1-��7L�q�5*;??�:%�uF�c�~���F�t�l�ʽ[d�?����)�~�̙�A��_��dמ*��'��8Z�N*W^��,zl�L��{%�N7kX�]@�ؚ�BY��������՗�nvqCc�46���3H#?�l�����e��"�}kP��Ƹ�V�;NO�d�+��;gȌ�#���IWs�ޯ�k�3S���'ɱS�ɅW>*k�H�Cg^e�+7��P9�}5V�}�,|d><�-�!!  
��+d͚5F�[�X�s�GV�p�\|Z/��w�HUu��`���x|�Kj�z��F����˟�8KN��aټ�e_g-��Y�>W�x��?#U���t����X��#�u�����o�>C�\����͑�+���#�}N�+e�[䞟-'��_��o��]R]� �����>SN��)5Mr�n�� W�����Ø
(F(EVku+FQ%2�V�u�r���l�XR*��U��g���푕,�Jk�fq��J�F��x����صߛ"���w�a���(ݱN�K>Tb|��Pb����݉�e��WL��zD���}^e�;�͑��r��ce��RIJ�Ib�W���o���
��/c
�ȅ����T&_pgTcֺoX�����m�H�ٴy�"����2u\OeK�RS�h��#E�o.uv���2E\��x�����c&��?,������
"�UVP��C9�l雗��v�Ab,ئ�n0��:i�yґ����[~��RY�M���z�{?}O������ҝ�7r#A�aR������Fe��N%��H��
�%�>?�(�����!��&+9';IW\�Aۿx_���K���{fF���U[H���2�G��f)��kŋA~Y�Ab4b;i�A ��/WeZ�N�8:b��F���)���Fz�<��&��Z�+��jw��8�i^��=UR_]*��i��ϙ ����M ��� i�	RV^�ȑ}5F{q�0��y؆�����o�x���vC�r�Ttb����j�So�[O�Yţ�L"R�qd�e���wX��7G�����;�c�9
�)��l�X��I��'����d�`w�d%Ii�#GXٰ��D'�V]S/{�5J^f�!�X���Ȗ�k���#���Ęf���� nϾ��̍�@�y�{J�^�r��CU��5;ο�@�����/��+�T�iI�Ĕ���q�All!�66�	՞�gw�1I>x�ߊ�:=��	#G6nq��p��~=�)�͖��G��[�ad�{�)QJ���I ��d�V�]�!���n�2/ZV������K/�dvq��18��6�\� �3D�y��ﭒг@R�bz�;
����	a�92HTb,̶vJ��Qr󏐵��ǞY&W\|LP�쑝���k8���T�?�}�����'�EU{q`�6N>xs������q�!�8v�@e��Ab����:o�ߒ�䌨;�Y-�AGΔyy@ޝ�Q��rQ[�<Σ�q!�3���(�W-��!3���"Db�˗/7n�~���D���G��)SU��N���~�%2lH��x�H��X}i��F+���*O@�Ϳ{M���i��g�Dod�^ϼ�N�_y��K%;;U���V�-I�NB�x#7�r۽o��M�2튋̼�1��<4���W����z�����a����Ӣ��IP���R��$�3j�s�q�ع�M��(";��w�5���1��s&ʇ�+T�M�|�=�6�䆟ɏ��K.��x饚;���o�+�z|���6K&�^�lV�k�1o�ae�)�����1�R~z�q�B���ei��?�#/,�Ȥ���80ٹ� kښ�"9���W�LQ��@������a���r������t�/��q0�]��u�WO��ɓMX�
�j����c�k�-�!~��������-?��L84K�A��(��={kdgY�d�<U�~�ʪ҃H3<<�^�g��e�A�O7���]��'d☞2����k���5����5����Hbz�Qm-X~�
�_���~ ;�����O�}p�Y�#�z�� o�U�e���s��e��s���B��!����6�*�.���a y���c.�����TVmZ!�%�ū�+}�9jȑ���� ݽ��i$e����Kzn~б螷��{����-�d�ƥ�֢�FcJ�/��3ɸ��m��H� �9Vr��s6�K�C����Stޕ�p�j�_W">�aه��)�����&\p���I��w�.��]Ch���hH��5o��o��0ZZu�f��p�sN�d�%�.��1��*蝘�Gz���~BH�ə72rɽ�:QrG��6GecD<�1gވ��y�b�~��!8q���®`G����x���!?D�TĘת�!;"rq�o�і� �yc�3os(��ɶ�����,Q�z<z=o������jYhP�����/���Ӎ�E�	~~��a)R�v���E����(q���^��� �|w`�d6R'h�[�*B�6�9������!>���3���o���  y֬Y&I�"DCT_~?��3C��_~�e�k|q-��{���>������<���Ki�A�cSe���ciA�x�bg��xꩧ��N$�p�Q��裏9�q�Fy�wė é�hb��8
C��;��c���ůApjR���7K�����p��/�ɲ���D;�7E�Q����^��J|j�7�oSF��!}����/�-/�چ��d�z%��(M���)��֔G8;էc=��c�H}S�|��"b��_r��Y�I	q��Ty|~��'5(�N>"KR������A���2���*�|��s{��Kf�7��U�9���	y\����Izr�؊Z���b|��+���D<u|�Y��,,1�fGI���N��u;k�9A�"�oR|����OvD�����+.�
�A���� ���Y�Z!ߜ��hۊ��Uef�����Se���^�j`�D�')�����^6�3��=vH�D��mv��\T/[����2@L�Щ���;����ʥN�N��}�y�N��t���Qį�V#��$^��6��������17��=L���k+�̱p��),k�:�����|y��r���ʱ�3ewY�4�[��D�����d����g�HB��7.5|�-Z-�,t2�T-���|;fJ��i�qf�r:�Z�1��}�RX��K@liu���b䎹%R]��w�V P ���c!pM��KG�׉���qeO�yڮ7d��-�+�T:�_���JaSd��dx^�<��^5�[�`��v��� �����)HX��u;k���c9A��� ����<�v,�\e��x���;K䝏ˍV��/'�9�^�Wf�a[EM�k_���%�D�n�wV���"�Kuek�(c�`��݂��sXЁ���,�3�$O�VR٨�ϰ"V��χ�~����nWM�N��0&S��y�҈�rK���ݶeo��M���f�F�o�,��Ň���O4i�6ށ7��؃0�X �6,-
�@�HeQ�Zv�a"��.�!�Peez$H�Z�ŕM��R)�j�0 ;��:/,n��}q�>٧c㾌;_u��=�g0ySii2x�`ٽk�,��m�)�ѠN5��gL�8o�*�^_Q�\H��=��A��פ��}a�HGE.���ms��	b�ymy�!x[c�X춋��Dbˬ}�D�����t��ҩ ??_vn�&K� �A�u��1��'�Hz�7��dm�]'��WF�q���c᰽c�
 E�,t�
b�]�z�!�������-Y�dI����s�1��t<QE���铝 /-��� PO�'G������w�����~wbY�<�B��p��4�����	��������5t�Eň#�����)�h4��?hA��x���Z�I���Q���F�N����ފ�#GP�H��[��t��T*�\x�&�Ǉ�E���_��C�Ô��q��E���)=Ϳ�T~���)Ƶ�9 �;i��4)S�m�����~���:*C��
� ���Ͱ+`Q�k�_z�%�e!�����,N��ɥ�^z�����T?��F����k+Je�jZ�(˸ٱ�Z� ���6��țE�dD�d�^�a,��D˲�������׾&�<�1;(4� �Un �$\�_ a�wךh��w�E슺�f��o6!QU��d�aCᮓ�6W��?�Q#���F�ފƮ���$�m�ԩ&Q���g�}V^{�5C�0�C�������8bH�	}���Mmz����V�I��ũI>��iʆ>X[a��l6Ao5 14�-J/��U[��;�m��� �J�޽{��ˍ>����4�>EV{�]���o\'9i�&"�Ya����A�a��_W;y��FTq°tc��7u���� {�Du����!�	'�`�`v�]�$p�� <���{�VY�&h�oeC�BeƤ�Fi@y���ii�.��B Mz �%�<�Z�*�P_A��A�����e��bΕ�P���������p0Z/o�ʛ[��<��kd���6Y9�,�E� w��/� 6 ��&���o��8Ot�kdA�,�Tm*sd��4)��aCh^�J5�c;'�Xe�ʭ5]j��b$U�Р��H
.{�A�zx��ϝ �bx^rH�Y�\�E��l��=tGʝ�4�U6D���I_௯,�)�g��66ICWʐ@�������3�qKM��?�|���,+V�~G�xx�	D��xB��q�/�P)o�Ժ�]��į�@Ö�u2�"��+��x;�z�+wrb�a���W\a�	���'��~��"�����J ka�s�8n���W��eJ�W��H�����yb?V�w��&��������#yJ�:��r�9Bl�8�!h�C�&|�nۮ��pH��SO=%4�a�!*A@.>({�UWy\�=�9�m1(��x+�A-�uҨ���+6ε�a/GI3�E8��8ix��O6A�-E��dO�!R4�C�����VXTѵZ��#���$^d	�N�������V�ߜ�D3f�0:5�0J�8�7��_C$W>/����T�;4Sm�����Ę�qy��p�z�if�%H�� d�'7���:�Ⱦ�f��ۘ�߻:/�P]�~�_�n|Ʊ.�&x��G���r�6Y`�jS����G�L�/5����$&����� KA��1z�"-Z�
G��;��T%J/բrt�3_a�"sW����~9�2�_����u4v����+��X�:;�o߾f�����i��v�te��5��v��`V�*\�XIZ�Wv�8�`&K��Dg<�jXRhB?4U�	�l��7���j��
l/i0�t蛪��jv��Bm���׿6��/���}�٦0�̰�o��4}��H9bB]���#z��o��b�X�P� b[F���S�e��Ϫ�C)D�<�'K�&��OV{�n�z��ޙ	����bR�
.uv��nM��I�g��|C��j�W���Թج���׿�e���v�i��B���QG%O?�t�	`���`U�$�b4͇��Ak�l��3X��d��&_������l�ߐr��#6E�Ly�G6=�N���~]�]�Kl�&�Yw��	P��!�C5��&b2ā�ݸ���y.���Ξ���,Аȟ��C,��!ҕ�Z�Y��C|n�CM��RGf��6� 	v�8���Ů�,rT[3Z���O����t�R�ԅ%�ǧB�v�DC 8qb����:a��r���,-�=�fţ1���0��`m�0��cL��d��GC(�� ��"�q���թ@�8G�?���r�uי������T/êº:�C��
���O7�%���af{���`2d @T�'�1dՃ�}��mU����O�el7ۢ�g��tY��p[���SM���|`ކ�]bm�zWc��b��`:��7�鮩�
���������m>.+�,D��hP�T��)kPA�J��v���#�EL�ú�dk�ݠ���[���v�,��+�m�(+((0JS�XY��ّ������{g���a'~Za�%���U[�=���j#kI�ț��V�1��p�WWB�l�r�{�����$�6�j����Im�u�=XS��E�z�hCMK�aSM��C��@�	lu׉���k��ӛ����x=��=jQ7 ��x:�[w�6_yp(Z1��	p4v�mj6�W�.��'O7V�b�I|q_"�'�����&>`,�i�B���iӦ���~!KȘ�-f����9�,�]���h���� ���y�xĿE˒�������w<넁8��w		t��w6��-�Ƹl�m-+���&����T�v,��]��] -�^cx��e����i4�g�ظ0��}&?����,�lMp�E�����F�W>�L�vZ��΅��.M�ˌ�n�y���Hqe��+�ND��c�>����}Yx<��ᮤP�`����m�56BC�dkjM]`�4L���� ;X�''���J\�<�JEVzs��ek�]���B���D7�K!$���3�L�O"�c��H�ƽ�lm'#q��d�*��,ͱ�!�7,����	�9pRw�pX<oر�.�}�!dH@&�w���z<�|�ȅwה�5Y�!������RS��a���\��0�.�<ei����.�/9o��K�/�$�{�P���4&x�ǂV:�!G�H{Ƣq��.!��{m�_�I!� i�x{�����n��p��`�I�t������ԟ�����$�ט�	�o��¿��`ߤ�m�����E�Ŝn$�PI�h�Ð���%)�qR�
PA(\�+�և8'�H0;���$�C�~xW!���2d.B��¶b�V !|�&E��>�������� ��XI�����C�����o����>:S�\P,q.����lA�Ӄ7��X�ZSx,�R�w�{�9I��V�Ww�#�����BXԨ�,z
v�$��w�$������]l�F1l��-D��LS�X�Dd�2'V���Ǫ�k��;k����'c��I<c�;������~�9D���5�6w��Pv &y衇̿�Xz4���<�yYT6��Wl�1�8�:t�|[92� C�ߴ�0v��Ϧ�'Ȋ���M.�g���Tn:�B��?&~ī��P/��îx����N�,`[!�݀��7��w)E����1�4P�+?2E`{q��V�k:9d�U�_[Q�dǻ�b��|-�f$�� �S�F>�Ġ����f��զdAc�˟e�� mX^��d�����.&��O����|o�Q�ρƌ-S���QwESk��n�#C'���Z2≭�0B�o� �$����k�4��x��w�I�c�G��`�;���R��-m��Ml�D��_�u���pv��:+�DY��
���"���h��:��v����������� ��u[�P��@nG�u%X�XW;�ŉ��x��fnl=_[t�=�6���l�. ��8a���Z�C�䴁g<�wSM���l#zsP΋��`�0L@*�M"�z��
2
Wms�O|����A�;���
r�P� �]���%���	V;�(^V�0L[�X���ɟ��'�$G˾�
����o6�YQ���j]�:����,蟓h�������^|e�-�}g��dD_��Ѝ�������JJ�z�}YV��\d�8��sx.��7��Ұ����~����\�gN�a�uV�W�\]n¸Ѻ_��N�|����f{M���;&��,V?�E����vc!���j7Q�=�����o�&y�^(AL��D�)�yn��R�~��=eцJY��ڴw�uB�W��Ū�� �WB㯊�%`��*~9���i��<�m�s��`S�_~�! �qd,��?��pm)V8ķ�e�9O����������:"K�_W�+��$���J0)A�+�X	QB�`�B�:*9���f�,��)��b�R����#�Mׇ�n�[��|�?��O�;��E(�`q������t�����R��g���cOd�����،Z���C6�ݽ��=TV-W[�*��}��D6;��d/Z-�*?�<0<� ����;T~yzaI���_Hn�(�nvRLA6V=����-���AHV<,���u��֭w5X_�o� ��c�1,ş��e�������'�:�EJY�J:��^��Vk�(M6�G��B�2��S"���� �2L���r8lZ~�.���~� �����w�qH>/� Ų6��|��̙3M�
q���7&?�	7�tSTyb�NrA/,�ՂgFXP�s��qJ����%��#�#�ߑT�����Gf�U�+�7Jr�	(I��%��v���!;�`�P�ЮP����?���L�ܝJ�*Lw���p iu�4bqr�DZ�-`y�[�a�õO8,���+��-��>IF��;�p'Ũ;hXoji0���x��z������`Kz����TиPy	\a�>�q(�/�����ch�A	 ��Z�D;��aD.q�ʭ����h0�!ׅ��?���^{�r���{┅�G40�l#�V�uCa����E@��� ��|�»#E4����
{��z�3�zDT�L���J2(�z���`;`��4�[*r��⻂�c���M��n��CU���8�Bk$����b^��:���z�T��[a� ��L�	�/:Б�� ��K%p��!+��HU�_��2 ��!q�����u�����!��C���i)��w�)�AI��\�3I�q�v���I�&9��h2W
�;݃�CwH�dAr=2��*$X��U`;ʡY��G�>��!������ �d~����"��[Kq���x:�Vo4)�MF�#�Q�I���=g��4+�a\���z
�J��(�tw�sw����fL�PB��G�駟JqQ���^'�a�+�Z��m����~6!��+`��+���o;;�]A(�gzp)���np�Y�29܆; �0)u#���P��kdO�Y��Y��*�b��7A��7�4�����r2����<]3cL���-�����o�����M2�n(sx�����3UgD�#A��X�$~�Z��H�:ݼ�1�0�L���	�$����.uH�)vH��5F���D9�= ٰ)� ���ļ�n1l� ��d3����߲i���47��Vt��c���pD҈�ҍU!Z�7Д̨�^'N�)*k0��`��w֔��v��N���v�!m�	�����闕�0Dj[��rt���;�=���pʑٲdcU�1\ t����-��&Y�&�3_W�+ٚ�E�(ma��6iҤ��B��
� =)@ H�0����n4��`Y�nք���&;�E�����O���Nt�O�"�.�	fB��K�`��IT2���w^0Sc���t��t��-�u��K�J�k�"�	E�g�u�>$<��Nkw֚RU��!Ć@Se�T ��^�:�N���;��|�ȁ4l�R����f�qh�x�E���1/z�V����ɼ4� �V���0�9�͜��e1���6x�(c75���cu��7E��B��9�F�H�!�$<P�jGյ��!���n���������=���Bڏ�3�˻���\[~C�u�RW�}Rp�p0;{�ؘ���i�iJ��h�!��.`�3�kk	��t������ç����������?Op�G�6�ڲ�X8�E;��S�ۉy��sQB;�� ��[�����ilj}��RR�Ȥy�����벮d����Om�\[��VbFgǒ�F��X��JQ��,"�L|�qm!x5�$�KCRRR�^�DO�T����'��r0��Ma���w�3�y��k�KQѮ�;����l3v��n�3����W_-Y�Y��ܹQ�Hj=�~�"��?�P��|�56+;K.��"s?�T�_�|��m������7�a�<l��n��D���Jq�[O����9��2���*[\ �b�)E�DxVO*ՁiJ�F�y[NN�T��Ew&�JZZ�uw-�7��ǻ�yw�;��n������ӷ��y�Y&��M����7jēE2$?_�y�9���/͑x �X[�y�̙m�Yބ��hԿoU�?���[%*�&8����Y`�w�!+����(׭7K,vɐz=�Dmm�|ec�&L��OG��A$�G�p��	�| cC�h�� ����x�� I��v|B|̱�L<)QbE��=

Z����>�r�s����}uʔ)�_}�U�k���)���AN�Ȉ�
�ڮ\�T}� ���Z�J<F�]x���|9!�r@q�/E~�4ü뮻�:]W�lYү_�Dr|6�DiP�<r��1 ��C�@S��J�B�)}��:P��ލ��ڇI7��~o��������L|^c�������<�a��(Q�Z�飼����u>��]��������q���j%H���>��?m�,��񇑛d���J�A,��:.-���uXEQm�@�䣧���i~Z����t��ȓ�L��4�o���L6M4��L=�p
�yْ%R��H��k(!�B zø���j��`���^�'e��z�=d-���%�j9<i.] �c��c��l��p��ז:p�v�9�����c��Y�<(7��"[�6\z��6oR�۲cG�Z�>b����a��ٺO��k
��L"GF�3��5k�.��8����}�ň7|���6x����{�rsH �M��U��'�b �?$d��(��\��O"{���N��'�"��߼�̂bAd�� D��o�86(�����bR�k3H���hK<0	h������f{�M����L����?_����h�����s衇>AT�7I�<�0D��曏�gK�(Rv��:CU����SSS_��� ��I�2o#��DA4��JҘ��~���7�
�A@������a�}�"�.�}B���� =B�O���l�~b�7�t��7��A�%��6���x.�3�-[��3f܊������.**���c��`^;��IЭ��^��:�c�٣ǲ�s����۷oϡg ڃ�E &q1�R�~�l��ްo�D�Õ�g�,�Y�f�����E�O�0��)�'�	�#��Bj/���XA^��:���[шY�j] ��g�x�\�E�\嘚�(q�����ڍ��T�w�����>~�a�����n�՝oP��	�:0U���"���^��ICYE��lKX�;c�>����<^[ K�=���3�!|�q���ܰ.x0Z	�x�qӥo�L�x�֭�`ڥ߻\�u~��{�9�d5����e�`��W]e
1�O�S2��P&M�l�s����:|�OԶI�{O5����ȸ�ɾ��ED���1c��{�>37����S����N,Q�fԇ��6���@�=	�S��֣U,l��`_��
?묳̃�7�Y՚�.�f��#��;��ew.fơM��Z4��-��m�b�y�7�P&Ƽ mlm��a_[�w��X����^����� G��>3�S�e=��S�>m!Da�^�ν�xFp�BR�'!�8»U��X�p�Lȃ�'uoyV%+���ʰ�`�Æh�ikYm�$n��p  �@2Id��؍n���Jq$���������ޛe��ܯ
�q����]�=Hp�柬~[�a�"c1��n$�k�FN� A6���^�wV��31��@�� '�m��9��]�| ��j��f���ժ�zN���w7����hv�U�16>p�B��&��}^o`�/0v�~�u���h8툽��� �u�嚶ȳoR�����[�B�t�uy�1ʧ����Tu��3Ϥ�؏^|�ŧ��8�t�6�f���c���o��\��+���cC
�u���=��L��e:�P�|��7����M��`��f$�8�U��� ���3�x���u�H��={v��D!�x��Ǔ ���ĩ����(!c�{T=�V��y%z���_�W�}г�}W�ࢋ.�")Ĺ�+ڃ&���UbD�E0G���� �`�灻/��_A��A�|E�n_���W�f�A�|E�n_����[�V�Ax    IEND�B`�PK   '6XR�\"# � /   images/16f29068-8fa2-43fd-94bb-aa3b1aab738c.png�|eXU���B��Hl�"���H��Ҩ("ݢ4H7X` ()ݠ�ԢA�.�\�t�4��Xx��>��o���9<g;Y�9���1Ƙ��/+AJ|����J޽� �9����m{�\�y����-Iţ��zT�5����]5���&�0VT��ԶwTm,lt��1���6�u-��-����`0�0��o*:���l��b���/������q���<?J|��yV]"l�G��ׇ��?�8\���ʹ�>��N��p�+�{�+�=�������_�~����R�sK��0hb$��������!]�\��|1�����q���q�.I?�_�~�L𿯕�pZ��E��G���;f������!
�|���X|��`y�<"����F>�������j��Tv�q���FD�=t�{�\˸U-��k�V�NF+p��G�ڗ�+]�(Ǵ�=���}%��|�tB��I
~9O��K�\Nc�u�������}�������\O�D�[��oԖ�����
����}Hs�ş��r��8�\W�4�DUTT�$�ns�nľjܑ�����{��b�i�:0g?�cձ<V?f_�fr0C�U��q�+Q\�~;
�c�#"]�%�[��6�N5�]���^֥2��e�(�%�w����{:�{0��՟b��X�Jh���v���Tj:"�pn�G�=�`�?h����M5��AÇ�a��.�ka���i�_}����4�*���硗y�%�ڹ�m�e�T���S�99<�cS�0+̼Pre�Q��r�:�:��V��R��\�~�i�`�KE��Zƙ�t�^d�n<����9�﫩�����x��Z��?u���.q�J�<��O�C��~0����1���vk���I�q(Yih)`7ߑ���S��cf���{�/�n����Ɇ;� ŋ�������M[����ϲ��r�Vʨ�4b���9`x�G�>|8bʹ/�8·Vp�����T�]���G�]��VK����rT�:,������m�i�;t�(q^k}K��DZ�os��X#|���c�fL���YF�;�,�rg�DN�d���zz�	�����_t����?6����x���kf����^�r���oTЇ~Vj[^��&2X���������I��2��!JJ~��gW�v���v�3�Jì,���y��%�K�g�&)�����X�R�o��� H���)�@��E�E�8�~��HKZ���*萞�����l49�!��yRN(F-�`�Sfjj��{��=�U��|-?��ϼ���րo�.�m�|�1^��r�4kf������t��7�\�9~��)WY�j�(�l��1�����w����;�q �`�q9�Sz̤/.>~��u�FX@�w�QJ�$>t��7��".˄�ّ:��I���1�m_��.}s�QS[ے�_����.�U%��QO��7��#��.Z�~]�͐�Z��_�^*F�g�;��O2Z����UWDE-��֎���O��|�Jj��2��}[&�ʩ1?T�?�ՠ�E�}�'�\Ŕ�m���5J���4�6�xJJy��]��z���A߾��uPq:'�(��f{�Q����n�������j���&-(���w�{��VJR�YH\��CE'��q�#�%ڲ�>t�;V���4�c<<N~)�bґ�DLJ����Vo�M�̼O�U1͜y7Z�k�f����	��}5�{���t�>Œa1X��h�VQ������h"�`m�/��ā�yb������]���Q���8���V#.�Xz�Y�i�y�~�*�`��f>���B[9�(뇰��{A�M����P���gy\N��&I1���2�~�R�?Rv��.�λ�jZ��C8u����lK�E#�!������3���D��sɁ,*̬�h7����젦u���ʥ� ��?��a�����]�g�N2ʶ�l�����6�fp:�Q�:Uc02���p���j���"��������ǔ�n�|���v����o����s���+׮u/_p�o3�#Ͱ��D{O+�������^���]?�P�Lll��K���z���Z%��3a�	��&��v<�)x�"b�԰�-��*���%Ǭ�*�y&J<�z�6�������qj��sv�B����P^� ff��tB���122�7�A�]��=���t���k�`�3MCIK뉔��]��� 6 �f���KHH�̃�����X�S!�K����]{�UHZ���c�D�b���`��<�mH�0 m�֡b:���U���3�K�$������_�8Ե_��1�@�8D�V5''�ߙ�e
m1n�}�����ҧ�����w�+���9ߙ�xո�0�����ry����l�B}0Gp�T���P�t�~7:�����S�6mfҰ� A��c��������"��&���55S���'�"G�f��M;S�mms���0����Gp' ���g8{Rղ���o5G
�t0����?*�G��_8�fa��W�ڟ���B��`8���}������k$�Q�A������ܩ�$n<|���
l���3�R�K�.�@:a���%�F����n�9��75YZZJ/u�J6�,�PTS3�ō�����L���з�ii�l_*���Ƭy&��h�d���I����<�נ�jwo�[H�D8�;�~��K&JD�Ν;R���j�F.���x��F��s�>�N3+)*�j~o��x=L�Կ$�C�\]�殜\�m�������z�I�y���!�֗�0�س��^��@��F����
����]�2���܃��r=>Rq����̡�������C�=9�g���<h0,��j6�_���ryZh�T����l��H���jzw3)m0���cR�^�
�#�x���?(��c0^(9#�V�����P�&�������9����.�^|#dvk�G;|�����?,��r��K���$�X��͸��ı�i�~I�7n�3:3�]��~��[�áQ\�u�p�}O�|�ΝW�!qk3]a~�?~�<���#q��$�.<�D0�����T�繞�FK�*� +�|�J"��o�(�H=1DLIE�~�1��:�P�l��+�[��8p��T���h����G�W�3^4�#x��YS�Ы�����[k�%t��Al��iOVbi孟>�G�;�Ȏ�z�C��2���͉�.pv�����vS��s�.���Zmsl�.�g@e~���oQ#y�B��4��C;��D*�(�E���!$d�E�?IgBogci�5�]��鵑�V#U!AS�#��J�#�����J�ZԐ$m4A-�@A�-�X�k/�ˉ��<v2�q��� y=M��c� wp������DUs�F�O���NLL�wgϣ�o`U-�/y��{s�qz�}�%.�_v
E�7h�&s�B��J~���A׸c'/Or�oދ�nmmͱ�SG��4�^4�@Q�}Q8�z.E9���ʥ�i��:u���ԵI�>ϓ^��!Q*Ϙ���{e[��$/�w@� G����F�����J�'���(/�6T�>��75� ��S���M�BР��@RY����U��{io�B�ܽ`v�'���k&
�.��q�&У�"�&'ZA���
::s)��=��/�#�(�c�C%[�kE�mW	�����˒�~�/Z�����Pq�g�u=�A�>�1ϘXr���9MD�:�(*C��`?��xQ"H��cAAAVOC6U=W
�*C==����?�ܵ�K�ҹ��М���쑯}s`�߿�r(��@AW7Fܗ�9@,�(�X��1=��0����sXSpQ��G~��zi���Ʉ]����T�E��'PY]�N��(ϵ�u��mU-�˪en���h�`N#�����������˗5S��||�7o���K�X��ӣ�$�@aqw�S7\D�f�>Jd.3/��j���2����hJr���J�N��k,�%T�)i�]��~v�-T�ɏ�'��[ ?H��g��o������:M@M�|�y=!�J��x��T��3�Q6��p�۵��&�k���&�N`!��]�b'`=��)�(+H����}�������Yp��A���|E��;'	��
߆7.�m*�X�{[��[/ʞ?ޔ�-����"Ք�y/D�<U^=�_���.2�N�5��W������EK�s&!!���ᷯ_߿{�f�hr���&%%ErmrJ���|��5�>%6����>�y�s�PO?m��P4��/h�f&�]�n�p.^!��� H綡`����ի9P8Ǒ�;���E�jv�{`�L�Z��K*��J
�����m��.�C��l���R2J��n��<<���2�zd���:�(�>��#H@�q�ę�B�EWxxV�	�-9*ji=�������fm߶�JX|�С��{��xn�.e=��.�	7�q�Մ��qbe�����䅯$�r�p���jߙ��f6���4@���}�N�,�����*�������ՓѪvЭ�� HH���L�3��\�|꧑��ngj��AK �Sm�TUNc�ɀ̭�8_i�C�$b�(9:�T��Vյ�HW���յ��9�/rX0 O�H���yii�ظ89�-���� ]*��S�
�Et��r��NNuuu�;V��Н��T��:`K�D7��'�N��_af�����������$���i`Ev��}O��J��U���M�z�8�|�R+������?�`�Tmb����y���O��y"�P@���=���q�^kW����ȭ����Z{3-�!`l�� 6��0
���ϾH���Ť%�r��EZ���L��I�SK�G�~Q��P~i+�jq��<F��m�Ӓ���.���n}�����:k�w��K��h���9A$XYYY�@�üt� �� �7u�-e�f�V�	f|uVRR:�sS��$瀼i���YT�ǎ#�s�i~�F�Wto�E8�/aw�*åKW�����s>�̱�A*��`H���M5��iE�vV�˟��U]N�x��Kn���W�ѣ�_�~9>4?7^IHL��311��Xn#���Ҋ�e�!ۑ>�ټ�|U�"zs����&G|E;�sD3F:ޚ��Z�\�㷎�N�
s[/�2��nٖ��q/	b�HLMM=�t�%N"�3�� 
��7��W'!�E4��\��:-%`�vM��ׯu55�G䍍��ы�nť�6L��W#YO�8p*!>ŵ��i)��a��J)ʐ�/}IO�_U2!"����q5+�f���n&�4�@�l�����fuBt�g�Xd*̢����W�����~x�(x'�_��)�le{#�W,a�e"��P1�>q�i�E�i����C�~�CCC�����T�~ǯ׈�\�rWRRRJRR�����ve��<�����H ���ji���*q�m;����X8��营!36�磣z�������s�����an�9�5K�����,R��|�ʞ��3ok�@Ґ�6��Ӽo�@l���].�d�V��1�'Ca}��gD�_�m=�]��-v�����}Sg�p�։'��䂫GZ`�@�Eh�,o �i�	2�a���/O�/�I���*8S�_.���b֚��J�s,q�����?9�=S3fm������40@?��	�e'|K�}�w� q���OM#KF�[k[�)9�S�QBw�W��3>}Dp�j����g�������Af��T��?PP�(�3-�dOav�Խ""�����-�H�����6��������I����h@}+_D�1<5/����e����Z]N!�.�/0i�N��u��I��L��!|vQ�}o%��3��_�E	�I&`���=0�hɒ��"�"���M'={�ғw�~[	YPdd:�B�x�DC��F�ְ��Iroޓ��8�� /��
�
N��0�)@.��^	@����Ȕg:�:PW�z��>od�k't�i\G��:P⢤���N�"�֡�k7����Ғ���ƻ�#8�9װ��)r"��	��<��Q���y�J:�c6X�%�E&��t���+���,f�ܷ�܀^�W�h~�׊vMd�O�Ҧ�=�L�dg��r��TI\��^�����\�^HKރ#���k�#�5n�/��J2��[��K�(ݒ""��y�&�a�I�}{LG����ߚ����;��:ۓ-SK�z�h��)�w���t�Q�)��"{��\�rC��M��`��ЕJ����,���l칡|Mv��6��������߿����ݻ�����%�_YE>)<i�hru��@C���9���W�˗/�,,m*:O+_\>1F�)~��J�h��� z�1�����������R�r�zp�t��DS�Lmc]]+����f�'��H�YBJ6�JGA��W#k��gG6�	m�B��<;Ƽ~����w{}�[d�LG�C��\�]�������"�E��A��G��_?Uu��^�	���D�u���0�V��eJ(�� !�:[����0�G��o��QIЌ{h��vGǐ!L�D��m2����!�~,����R���[(?Em�t�ҍ[����a�::��g���YT�����'�?}�B��O�r���8{H��K{�:�ŋb [�ȶ�v�- p�����7Z	����ʆ�����;z�;e� ��"��{r�Y�j=-���rZ�w��	II)`���h����%'WY��u$ܣ���7�J�T�J9!�g�9Xb#[es�t���d����A�<��FO��U Q{�4�_��^�[}��}7aL�c*O�\��w�w����8IFV��W�жA��m=�˔�o^=��G�>;,��6�wJ���FC��c�@�6קyRY|�!:�
��/�{���X��l>���Gx��X"E������Q�+.6r(q~�L�Yf���55����s�l
Kz�-�W����E�Cq0���$b`�P�=���!ܚ�<��1C��g���8p�Z� ���@�[��2�o߽k+vZ�����߰
�fҖ(���=61�"�%�Z�Ձ���qE,h�Zj�$jz��(�t��n���lR\�"�'�����klT���-X&�I�����77gg�OAye5�<����t��%�kW����͏អ���T�~�V�|�x��a� �Z?G�|mH-��&)P�~E�vvs�J`�U��>����!��"ӡ�g���B�C�]]������R��/����vR-�v�y�,��7ڀɰY��G�5q�='%-̓�\�!� "l��SV��9JL�@Y���C8����?gx�>x�P?~<Sz7J�=���LD�1F�>�R���2h�|"u����,��2�A�SϷ�aB�����������CY3/���6��`�@FG������'���9�C������XQII_j t%�GI;~a �rJ��d033K�N�a3�mld�����IMe}O+�=�;�p	�- ��7ys/1"�6f�E�g?���׺T&��\qo�P5�K�~LK�� $��en%Lj��d�qQ����hT�jd4|�,ʟ����5j�����	�o�,מk���Mf0����K\�2�8�%��Y�AvO@H�`du<uU���Tp%�k �"�~�]&@��z`+���x�J<�L�(��Bq!O���Wh�`v��@F6� ��P��v ����㜖^��e[�.��xz"8s��OU����s��
�~R��:�ߜdL�̞���삁U�ˀ�09�y��x�kp���e�Iz6�Ǐ�0
�A��^)0��ǎ}-$c�QN��x����#���� ����HA��=�B@x�_ݴ �J98D�f��p�L�Y�'>q�m��HTw��Nh+��ŋ2����������ڧ��!��X1��lmk�5i��'D�yd~�,X?����
��zv���&[��h�z��Qqy`~�+��5d=�Y�$Y�ǟ�Y(�Yt�? ��V~��O��g�ނ������s�v��H��)�9y��я����V�d;ʻ�A`�FO�x_���P�7w���7����I��
�������dK��������>�w2꫷!��3C�!�{��&׳y��;t��a#gh���d��� �T�
T�Ϋ���Vd���U�v�`��M���8�Oc�e�0���9F��H��~���p�|���_$ �cN\�t��u�MT��_,8\fa�"�h�3�M�)�= ��[��`RC�����,����FJ0�M���壶q����6�4�8:�[[[�c-t�e}��ҫ٪@sz��ؒ����k�«Sm�`�ύ����>�^f�u���{������J��q�0��������ߪ���I���f����G�y�=�iU V�uݰ�{phO��ޠn�P�;米�����ʨ����%U�+a��
jHk~:UI���P�I¦]��\���>H3�Q���-�G���k^��4�zpR�l���,��ϿM�C�j_˾G������1�e7�ͥ��^8yA�}w��2v���1��B�j�x��� �n�2W���`���	��w3���G�C@@r�h�l�2��<�_P�X��qo�#�5����-�b��	�Ǐ�-9Jמu+.��z��|Q�S���Dә�z�(��l:��e`8�H�_aJ��� �YX���͛dBBj���-J7�=�ՓR���G�gB3VZ$���7^��F�"Ga�O�ѥ���l?|��q����	>�=6:��14����g����X�Jݰ���Fý��oN&��eT���"���<����T��^������P�% <�o}}�2u+�!g�%X��L�Q˭
OR��%L��D���/ᖡ� ���Ǿ!A�!��]��.&����8C��"h� 4��K5ݛ����oy�ud�"L��&��b<XZ�I�(�3n���L��)z~ j��4�$�c0 53��M3���P���������P�:uJ��E���ϟ᳌S	w٠8`�g�Duc�jZD�����̱)@݅�޲��N'ğ!�.qFҜճ1C���B�
E��`���7翼��\��_���~y�?c���[��#G�(����$�RS3mI���@7�`^ �������t)��̯�g��_�-pJ�����b%�~�C�A;H�v�1��<<ɾ�t*��0c�],Im�v�c�Ev�C���rssMMM�oȿ��B�p�g��F�����N��� ;²� ��o�+\��w�_�4���?���3���}���w��%v������ٷ8��t,W��4-������ū������L}��(L�}�w�O�kega/�����Yq��DD�8�IFY$=(-*�HB�+ڡtH��.wP����hjbR73=-���A���I�%%EPQE�� "��Okjɱ�S�u���G�����P��mY�y���R��'�S�ґÇ+���>EGG���8AGC3k]��}N����}0�(�;̍Am\E�Ӏχ�?{�'��Wr����2]jz����Bv\a�V����df.ܶ��v���������>n�ޅѫ�e`�61_3}���ZhP�X+:�U����{��x��4�9,S�i��%�}�E��?�:9���#{w��m���w�h]b$~/�1hdmaP%2�cG͹�]�����W���K���FQǔ�[��ڴ�;��t��0n�^���q��X������?�����ѝ���F�o U�\��@#�L�.��M2��ȼ��sn�z���+ܱI]}�o8�Ӕ��P_��n�0����qs�%;��c~מ�[y��c��d�i��\�Jܾ�s��uw�}}l_H�\�d�t�Ѓ�'��W9C;��f����3���le��L2�,� ��;���ԧ�D�C�Â��2�x���w;2��d�[{��,F�����;���ܼ�yw�nTέ4�,`5!�^��Spp������)�� �B�t�@14�Mӡ�!H������-$s;D���b��ݷ:`�������,�F��m����{��X�^���� v�Xv���w�ky�穋�R))*��,��� ?J�4p7_ad���3�U���o�B���M��Oה�� ۽o�+��V�(vٷ��-A��_##e��^�Tժ� (����>IKN�R���������!Ӡ1�_���ST�c-���?΃�c�*Y����\Ft���c�o�!F�*�#.]�G:	�тদ��. ����6��(���n��1����wo��n�����%&%������z�U����ӮÔ�� l�
����A�cA�����stt���Y7g����b��cs���Q���֡��w��W8j�޲�.x�2�l��ژx��eMII��ty�+)��<������� ����uzxj�ӥJ�(�.�W�������v{�7���F�a�E&�"B���,%�_�~}"���/��8�mf�u�{:�ï���/��d�)����)����/�����w����Ą\�5��Էo��A\tq,X�4�39����������J��X<�V�Б�=W���PX�Aו��n�τ��Lw���ef�
��ʆ�Ye�T�-//��φzROqqz���!l���P�7�ͱ\���<�~���|��MZ���Z�I��U�ߙMK� ��7�tf9�D�PQQ��F�y5���5p�7�e	L���VŬ;s�F҆�1���D�6����J}@�%�(?2^΋�vjXpрN&�f��݁?6���3G;��j����
ZA	f�:1f]�������o5:v�����Ԕ��5;�����Ҡ����o��ٜB��+W�|�$�u���/e�U�%z��������uy�  @V�C��C�!�:���"���>���-JM5���LS�P��\����olYZ�j|<���%:�VH)���~ѿq�m���U%�>��4��9�W9
�۳�Y=g�y�>q9�4^_�FD����\�͛ϴ��.����P���r_c%'	Z�CסTY="/))9�4R}�p��>@�h�+c?)������q0����4���5ݻ�����*b�v�,��٪�ie.�B��+�3�vA�.�9.�S,c����z�������傘�1�߼ys�R�����������8w���K@k��>��������*[�0�)z�t�Dlssen(S�[�f(��q���L�H�'�jZ�Ipo?!��"�Uo��E.JĤ//:������z��T���#͑.��~wC��S�+KY]]=!..nm��|WN.g޵�P�\��E��r	�ݭ7Ër`��f���j4��[]̸͓�`Q����(�/p钞��٬p({J��٤�/h�me�Q�q1/u�`Ӌ��r��Z�jkkѱ� v-t��K!����&ehR\���
t�g]φ?�)S~�b�4��rɰ�9���փ��s
�Ωc�q����/����S*���u�ʕ׏q�bK�l֚>��7M�y&(ݕ�D�3C����	���6������;3t���pD�=�,D�:SH��������ѣG���v�<NL�
ڋ�Uh�,���KIY9��iWz 5�t�#�-;�|Ok��?��>��(�r/>op\B��?{�<��{��0�в������}%-��]�v3o��_, v�l�	���p������|y��]Ni9�z�??�hҕ��I�j�N@pp��놯��>7�(ZU���L?�G�#��m�f��A-]����N�`Q�3H�=�:��;�4��>8f����99��^���,���� ߃a�P�N@(j6\��8IC�V�t������e�6�fZd�	P0x��$o��'mT`����\���GF!캅2ڔ�;D,aV�cll����ԗ��E$3�E�G�^����D���TR0?+3�>[����[��פ�0[�͘yO�����'իX'��חB�ļl�^!�2/���]��O��δɉ�am�Z/U͕��
�X蟮�t�����S�/����3����qp�FP�����z�c]``^~ND���@~IIA�[^��P���� Ad��5�k<]����,��)@}��z��	����10e�9Œ���� &���/ {ĝ��X&'�� ڍrv�DO����nՔ�t�����;��� ����g��l�p��ú��j�.@���DS���0�I/ "�����1����ƺ(ZI���mc8~h7���A���!�"��r�����&�����y��H��b��V���L�^��5���.1�l*^�E�7��NC��z{����������uttD�ʲ�3������+;<w�f޿�@���
�d:�!8���F:��'z�������瑂(���@�S%���*زO�C/ȫ�u�����7���-x�;(�⪙!��|O+b0?�@�߾{'S+u�^>�7W6F|g@ yX��e�y*���g�(~����U�VR�0�ֶ�DS�\��r���k�dŭ ���J����3���JBCϤ��%��tN�%ɕ���P�WVW��{@��-|�E�KA�6Ʌo���a�C�Б���� W�����y��}YY(>�B������ֶ��ly{��-�1%����e��EkP�鎔`<�tI*�/�t�WfTc��e!n�@Nf�n.G�wөFB�pD9O��Z���Y�n����1��=I�v洶xD�o���c�
-%� �v�����p$~�<ɕ�]. >n��@����$ڞQQS������-��M�ݓ�����G���G�/|~m�dY�Ul'�%m/�3��P����g�^����e��������A�p��Z���fҷ~K\�[��t)Qi����1Y�Jq�!\��jjЋ\��j=��R�ٹО���,����t�^��O��S�G��	7�=�e/ѝo�knk):� B���<��ě�������;ZZ�a(�mp��;;;���MZ	D"���Z�911Q�H��G�T�u�8����$kZ~;�%eR���C�<�w� ��U���C+��+�I��6����}��'%9�W������#�^�|�$	��r�'$T~�E�b�n���g9�B��1k�Κ��@gy�ؠ��"��������^��4l7��OL���W,"��J]7?�7����-�&|�q�nZq�;��CЙADD�	��ݻ?e��{�^�g{l:��M�v����/���SNU�z2X�4j��h�$~tt�uI
�>g0�Y�cR�Esy}� �gڟy���\%�C����;2�@ȱaBNY�ߏ�R֍,���ݻ�A���ж=�"��\`Ɣ���� �M������Q�m�/a�U!�6D
k<x� G�w��+p�o��뛛�U��:�,���ղ�&�);�D�7ߠ�8n���(�'G r�d�����u�2XpV���������f�^g�Z�=o
��g���(�	}D���*�9o��į��͑��]i�,<<�7wM��P.|B��0���Z�i�7�A��EcQ��z���z�/�"�TR�xAD��{���P�������޳�w�^�I�q7�	B3T�_9��W���#U���`��*�?[�Q�B��H�L�󭬷�g��6
ϋy�@���:+R�3�iݦ���d��;e�^�LCVMY��龿'!( p�s��Y
�"��^&�W05�Smǯ�������<�|{2\�0͞<�q�6(M�믗������m��GO2�z�k\�|���R�kJ���^4���L�6�_nm9�噅���nT��%R��m��_�_(^�t횲`��[翤��+��V[�v�?[gg��hN����*���� U�o޼�&� p����1g2���� ����j�C�+�����x�1��~��붒�����6_>�ݮ ���:V��M �,�	Y�NH^�o�9s��LЀڢ�R�uyy�G�>��� {�� 2�~�����B@/!��Ͳ}�N�����C:l����?e_T�f�}�őڂ�H� Бg��њ�Wmƥ���4Rv���Z�7{��sB�d��5�u����0����$QDz3�ٗ.^�T��:U�c�����f���|��[��?/Vc��;���*W��\�5hǫF��-�x9۰9hu�v.�������1�Yp�`f�S`�r�F�t�d�w����4������n��<F@eY���{�nD2���P=:66f�=wut|\DM]��y�Xr�����z�`º<�OS"r� ҳר�J�X�`�7�rVNS��v�����q���ύx��v}�^�ݺ��#�޾=��Y�����#st/�wƯ�"��� �EDD����㱟U埊���f�%pp���4
�6�U�ް��EF÷���,�_�d���T\\�{/��V������\�-�G�bB�%�I
a0KF,��=S��Yщ"���LvE������l�N��}�D���?�����ã#Z2�᫾�N�����)��20o?�e}^���T��mwj�_.��q���ꙓ^↑N�$���q�<<<9� ��EQ��sYiZE��@�M���L������LI��T������x��w�@�́�RC4�x5��-1d��c�pc?M��5���0Ғp!=��A!���|��OMc#��E�����nO��..//���5\R�h࿿��pm��z�p~#�e=:�ʽ%�H�(��������a����Eyyy�ʐr�ED��m����)���e����[�VUpr*H��6e����)�p�>G����G����0��>�]澟fڙZPg�%�u�����iPL;�:kR����X�Ms `a�ԽG���\Gs�dۚ&)�ݸFtE%U�ꖮ�n�=���lR�}O��H���#+���jٗ����� �����!���m,�l'�߲�kn�b:��	�1L4ci�1?��`��TH�Q�|��X�~pŰj�as������\����C���\n�7��~W�f2]��ZZN���C4ő��ݠ��!�]��\�LA��5�h���z� ��+ͱ��)	��_Y;L����8wL��[����VɫBb��0����2��v�WR��~�ldkn>/;wz��ԩS����:�_��E�q��U����r�M��az�Q����4��$+-%|h�����-�ZE�_�PPR�K���xٿk�י��K�^6�D� n�3���+��c&���� ����p�Ϋp�@�`hjH���ѻVVK[^�﫪v'�mg:�d��V�����b����L���WW�*K��;3�9�s$JJJ��ܦm�2�N��߃ۦ\�@0��R��7D#�>�X�#�O��c����ģ�>��8��w���E F ���)�O�5�@k_����{P�V�r-�//߂�)�Lc�� �x*��*S q�N-�D�ů_��2}�ԛ���}$b �Lll��YY���9�8�����0-II�����`T� |��?��F[$�)��;����8&"]����Ҧk���cG^x�:�'�R�h�"�xT���r����VVV������0���<DW��N_L���1N�H�Х&ɗ�"ă��ٕ�����PbP��q���������Jl����J���j����:�N����L[���{WJ����YiN��.�\a��,��`$����/00!B�sU��Ý;��^K���-s������%��&N\m#箛��=�mkJ7�]����`����}ѹ��w���;��[���$Q&,񀧦Z~Y���vg�.�����!�OȻ���U��-1�	Y٠��O�l�/�LDL���z%-��aK��!*���.���G�9W+�a�y��^��j���
ڧҸ�~���ى2Kw�]4�5%$_��+�IT�?N��a��Ĳ���-Cv>�7 x�ȿ#��(�e�r�k���0�.HӺ�Q�G�L���ₕ�^���6�'i�$^��~2 ��%4�ŜK�յ8ܮS￥������i���96?X�^1\�fN��u|��bt��J��N��k_�.Yh����dN+��I���k3��X�?��)ם�j���xA.r����0�j��:���#������t�Y<�>�I�:9x���fQ���ߏ1~:C8��E��~/��f�-��6�ϸC$/A�'�X���020��=��`n���W���$؂���珐�[�9�������M�/�
=B��ڂ$&���S0ؔ���$h?������y��m.?44����8�(-��\n�w0��rj^� {����ز����b�r4<��L`��":_�hܣ�K#�^�N�0o�:D����h�̻���	��vqw����Z�R���1|�h�&��#F�k �nV��k7'8�g� -)�
D����[?���j���?�|��\N[7ɰ}�S"2�Oc�FX�@f
ػ�g��w�Ɇ�V�?~�02����{V�=_�����H�l��O�_\� \-�Z~MB'ԍ�e�sY&3{)v��R�:�\A)�j>��3��1��<�`t�;BW
5�MNT���5�C@R��O�r��2��� ~����P���8B�^�GM{��7��b�uMMA�(��?�h6<��\�v&K�ٹ�U5���s�MNO�U��0Ud@��)*Q8�+��������8�n����]�
ۍv������Y�ٹ�>�]3�ʊ���N+��wM}�zۼk�U������U�nN|B9��˛e��\�&�>:1Q�o5B�q�|��߿�ҫ���Spgels"*x�Wt �� �yy|�F?�w���67�Y�Z�1�`�����ҿ|aR��7���§�6�r�[?��<+E1Q͔����ׯ���}1(v���s+l��&��7Bb/Y���8G:���$H��*�QA �6�:h�Q���Z��DG��@�<��&l0��Nˣ��f_!_�M4E�`	u>���Z��,���v��I��N�XC��j&^���������c�s�#U��:�	�ppX��r>󰯓�`����Zp��dt�v�.---��׀���+8�G�}E��f��mms��gҲ��.���]E�h8�ϯ�W�vS�����>�n�f�II�Ů���"��[vW�Ο�)X�Ce�A�ߪ�ؐ&Z�$��q��k���	>EI�A����cQ8X.���d���k�7v7
�<�A����:r�Z��Rm�TUݍB�[?��i�r�����n�΄l�DBii���p�?�P��0g
$�k��v`��4�ƌ~TW�3%Y�yrpэ�]Y�s��)bI�`Mq�To��k�����≍��,��-9���S��ILJ���D�Cy���w*�Nw�_��蒑���n�[�#����K�m�m_%o)���Cf�s����g��={{{���l9�kkj~6q>�_���m�!�� #�đ9�r)�qwj1G�h�țVPY����^���k�9eTsR��^�咯���,�4	jL
���g+E�ϋ��'�i|�ar��
J```�k��{:O����;šJ��HH���H=y�䎸xUA/����J���АE=R����g�YV#�sX%Z>So�,��`B���U`�r۷DP�@)����b ea'�	͞�g/����ROSY�?FS~�<�j�ǋ��`��(�h`X�YYg-4�4�Յzٞ�]��u?�������Z������ 6Ts�#~BҎ^��k��`)
�d���-��S������w �܊ �D0�cxћ����~�«�;�F
����ͅ���#�frg��`�.��h����	�W�)�8kr�����Y�"��S�tŴ�e}}}���F�h����l�{��(�U%k�,鐫w�(�u����ga������@2u�%
���9#'g�|��G�5��>�H5���s��z��-����}�F(���K<�@3���V,��廇�|)����Eq��!�c3�^�	F+J�"h3҆�&,W���%_PPp�E��d���eIu�Ѓ	@R쁼|L�W���Uq�e}U����l�������O���Eh�"<�V✋--����� ,���#�'�:'��-�zyz[#4F��7��jj�3!k��q�w��t��ud�Q�%�Σ����,��mfh�ze���L�bL�u�H�x�`޽{�&{��H�o�iF��|�d��t��b�F�0�����7��կ��\i&?��ٴϟ����y��64�ǉC�ހن��u��r�\?� ���sk�j��|��*���U�鉋�F0�?��hn��|ę��-z���(W��������8���ۨ��
�xD�k��r�5��bI���p�VD��t��>�7��لp6u�󔭶���g���  ,?g(��5��k�9W��t���5 ��.�����h\��D]v�YIɕ�s#�x�Yo��۲z����㓓���"� ��?"�eO�Y}�t]��խ��[�P�n�C/S����ٰ���?ޜ�0��5��_l}w<�o�����Rf
ɦ����2����ݱGˈ�dš���ǱJȖ������s�_������s��u}���~_�W�C��T�����r����w@]]���jǫ��'�P�^�zU��RSmՈ`�����]5���bb����?:�{���:Q)�]x�ߤ`ύ'�ѷ��E����{���MQ��-3��R�˅h����ʚ�S�#��E{�|o##����*��	�j{LL�����/��8z��lYf�i�ؗ�LĖۉl&zzCu�����9�k��PE�3�ˏ�ě�����1�7�J�D�'���P1���Zr���q3K�_�l3{#ZL��5�#�U�7����p�I��P��s1��n�����r4&�`QҞ����}���J5�!�-:�2�8N���;Q������ډ���iz�@��;b�ѷ��ĵ�p �;�bK�VrV,s��RZ��\�2�&I���=�t3�R}�yu81�P�U��1a7���=KbA�����q�d"����!�Oğ'�Q����N�M)^�ǹ�����\�ݺ	~��l���2M������`�5���ϯ8==}�̙���0������,�R��8��ɑR��E�i����ɶq�퟇PU!�t�`0<\%|��f��뭷��/����Rn7PM}�L��$y4��~��8?�����)��Ӄ�QW	�<��~�q���F�Ѭ�Q��h�0?�1��G�;���������e�v6ܷ?9W���
�<M��D�x|\�[7
g�E9�'8e�AѻTg3��΋+�s]Wq-�s���_|̷�'5�o���4.�@�%܅�oWёE ��o��y��ُq�BS��zz187� .� �xt�fg��ɱy��n].K�ZU�3�0h�l�܂����{!��۶@�����v/~B�G$|��莓Ԓ�,O]��T��'�� UUU5	�(�Ք�ɿi�[USs�����~a4�ald��Y&mk����H�A�D/��� ΀�{�w���FG�#��j#�C{��]EE=��t�9�S|�?�T�`�d$%��\c��/�%K���g����jH�s���T��ʿ<�c
��o��<	J��#g�'1L���Ǘ@R<�+��ۣ�:�vR�.���9;0��Q�dPL�@������'CCOݹ݊���,7E�̓ 
�	�t�/��';���U�
�\+m����1��� 0�[I�^Vf�mtB��Q���fI���x\fp^�hҕ-�-�̣q��a��}	����ܾ$$�gt��B�+���}�~��&IjK��O���]DV��e+���T����|����R��V��dh����
@���̢�TU��Y�N�?��M�"v����.7�1�;ުNX��	�z�u���vh��MKX��zb��T�ѻyꝧܴ���0@�Im��������@s;O�@Yw˅	8�B��5-#H>�N���(=~�d��x�
7Z��Rq���W��ޓ�d��I�
�L�����6�ZZ��J����ж�i(�Ҳ�޸*׼�����`ͷ���3�Zl/��sa0}��':�����|�����<T'����Ƅ�H�fg�M�U��/�s�u�v�\��/%a2�h�wo!,U���K�����N�����d6^��Y����="�hQ�81))�u����Z�J+F�e��D��R��z[5C�b�q�	�ޔ�y�1P���4���V�<����j�gPFg�)�C��~12���w���g��`�ǡ@�-^�o<�Q���`��-Ӟ*�ڳ3:;{��߼���y%%��Ô�#��������y`)�9989�6��Ov��><<<�������6������7��&�ѣY�h9�յ3���-O�4CZS35l�9�~Ag{Z����ל/�t�*0�nDfA�Ɇ�\�k(Z(��D���%���
`��:@of�m��iiw��
�y�@���A�h��|J��(C /������.ްis��)��6��j�`���l�2 ��>��S��Y��	�O���Op�3%_����3ȃ6x��Š4Ի6ic����)��0cׂ"��H���|��H��6�ѕ��vsZ.o~��O�J�,&U̐��$76>��쥤 ��.0p�ΏB��9Z�,��
s,�_J^>h�nk��X�R�>J��v5kml�����"�Z�Kx�����V���{���U/x(�Z(H)�L���/g�)�V�9����}0rc5 �V����+�qÇ���vӕ��u�$KܸQ�զ�bI��W|:~�<��b���L��!��
��kK1��w�^4���e���2 F�[|�ٱ'�F�"�+f���8d)J�궑�Af��u��d(p2O���{�r,X��Ҍ+�,D�r������gYXn���?S��s�q%5���)A��4Mb.A�'~���l�aܬ���c�8"Q�G))��P�x�n����?����<~��h�͵(-������a'^���.RAW� ��0|�/o<���$��e��1Y�0YM��v�4��t �������j��G���X111�n7�����bH�%���m�`a��b��Z-��ZZZV��#' N4@i��s�$_���w/�Z:zv�R�<��;)����h����;m�in~�[>X���)�"Opz:ߦ���T��0�')""B1���o�+��@��,,,�q=�==���UQ9/�!��tt����䦿�f�l�%�P?F����`h8���μ���!tFP݆�����ÊI$��~�B��ь_�E�FW�.�����ՕcƐ��R�*O~���W����� �,>��Bk���	YX̬w�P>5����
D���Zե&af��GV���!5+kN)���`^�6�B����lkd�AL� �X"�4��3��6`T0��S
�Z��"�j�����>��ǈ'�k����̪�����]]eS2�̬����=Ӷ�;��m~��'�O�а{zzn���<zt����������k�U�vN.���b�����?~��=�V�����:cRvvK�4�g�+�B� T���%oc}e�����-{�"x2��Pc�3�\�鑥�6�������8�[�4dQ��y}P������y NG�xzy�|�rÙ�-��n��M#X�:�a�&I7�-"��)>�i{m�
��Ž�s��v�X���G{t���cbc��_2F�F,2����$����:��hY/��ˬ��{�yfb���kc�EY��z!|]q��6�Ho:��=RP��|�NLf�]��yj���_Y���T�dF��G�"�&\j�ꊮb� ~�b��d\aDK��8ղ�d��z.UA���=�A?�^��!�_&�Ro���UCc����w�2op���W���6���`��ƌ���hP�_2	��N����-[�+�ٽ1�G{!����B2��~H�܁6פ��}����F��F���� }Y��k���������I2�_՚��Ϡs�EǄfC�H�.]ZS �L5��i����N��΃y~�Լ^ohd�(�μ��8Z`��q��hk{�oS���蛗.^T'�k�t���ǃ�_B	 7@��XH�b3����
wq�!|
��w�]tl�zʆʓ\Qjʪ��ム��s�0�����-�6.OT�'�F�<Zܺ���FRe���t�ƫD�6��Q8�]�s���`O�7G.�D�����**(����Ԡ��h?�]+~XB|��W�+@>�^�zE�>�������ղ�hj���6jsԔԙT��+!��`��Zk),�斖J9A�9�	�!�g<ԁ/���j_�ٳh~PޓZNN�roSU�n�	8`��}sN�u�$���9/ ����a����S�~����e~��'O�@1}
\E��:��u�0�xv�ӧO?�\�<�q
�S36NЋHL�e! ����O�"1P���5x���l��a���C�
�.�%�h�ϛ�ƻy�ƈ]t�iOAa���	^,�#�����Pd9�F��d�sƸ	jpMs�VJY�w���w\&�D����܊C�Cf����i8��	1W=������J��2!*(ǩS�6���Ѯta[&��{�<z!�p}$�f�2�u2	���]-�d�Q�BM��ty���ƞ�d�Q�IG�tSm��/�uh����{���B�F�Rd;�D��g4��Cq����ۯ�~�زH=1]��܁̣���W*�d*��6�@�2��B��W?�ĔE**��Kwf���{JJF�� ����S�T�lޤ�H���a����2�3�ˌi�̯`�M.^�T���a�	�8R܋F���T~��ſ|�Eq�`gI��ϯ��w屩WlTV��SO�B�
�Ɔ�y	���۷����Q�`�\��(c�:>t� 3G2����nNt{���g�p>���ie��R��ٔ�����C�~hKRV[U\��W�w����ԲM~ʧ�����;p��)Q��+!6�>|K-��$�4���p�C��{E�����ԧ�+����A��3:��������	[)��@��q���C`!��JH�2���J��ϫ嘶��xC��o*(F@Wt
5ut�!�eJ@\8�
�I�Mic�#d|�e��
������1���jNj9�AW0"jo�B'~�o ��ε �+)+/���1�����JC�W�յ���ڡ�[��A sM��94Y��BT���{��;�'z
�@klN&�NCE3�S�����[R�- VjG�	<%�e*�4x0�s|�?��5Y�f� �&(%��[���mX_TŤ>���E;��~�����(B{����;R�rccc���+��s�q��\��˲ 6o3���h::��8���������F ]\y~��M��:;��]��~����a�f�	4��@t��<��]i���fV�ښ�U_��8�7�%�$ ����ٕ+�SC��M�6��~�C�
Z+o�5_:aK�@d�5���(n���J�; &��(D{fMgn��'??�	@Hoz�M�ҳ��Pu�`/�K����A�Z�,� ���V�K��ŉ��^߷W�?~� �Ҿw�t���y���1_�Hc+�4S84�w�<iApr�S|�-��Hi9�78�b�A�)��2(lh����S��П�U�?;;��}+t<�"���
6��&����znn�;⛑��՜�"��3��b\�ZڴOR�w�����94b�%2�O��T1��H�yR�����P{�;���Tm6;0��ou{� 8��B���ء����ϟ��\z���72ϓ"���e+�E����/z�E�S��Dݼ��X���K+游D��-��B���@{�{w�"ǹ��6fm�[�ܡ	imD�x	��\�$d;/�[�7o��̇^t�`��X}�b�W:T���&#�D5677���\Ϋ�����lӰ�ɡ��Na����ϋo,����w"�b0L7�/�6\�l��|F�;Ӫm�F�^P�~d4��<�t^�/��.�����y�;����� ��?���dd�t��z�8��/��"eL�vv�G�M����a.4���8��K�:{��h�2�E��a�y�8�OE`�d�C:�rP_ܠS��i�p���x�����t��DD˼N�0�v����`�����@\J������Kˣ�8�ص�y�	���Jw$������Q`��L@;�YT�Q�nV�S<���\BZ�A�5�����	Hױ}��J�.�v9Z��h�؝���eq$�"�M�4Z���H�C
����`��$1}e��YYYfO��Y��d����[�~"����70)�K��-��N9�-ii�X���[��V��*FR־3�P���c��8�0�8hҤa
2� ��vW�0it�Z�����b�P������l�����ݝI�����Fe�v��|4�{+�0�c�^���C�^���̌�`>!������b�!���=���eB��ݻ�#���M:��}i�<C����f����+��P3s�����)�oK��\���_�/.&�¿�OP��o�<y���8S���N��zS]���j}���ҹG[��MC$)�?�.Zm�-�5�~c�W��-��U6��ɓ���7���b��P�Z����;���F*廎��O:3Go@Ē��[m�W,E��:k�|��1b�W���B�E�f��^Nw�p^��]gA���4�oA�������Jܒ�?A�0?�e�&�������������n���̌��늁�h���˨����������� �9
�@ȼG!�$$�mR�G�~����H+ �<����+j�U�,��
�A*���׃y#��:S���M	$�[rr-�5( �6��8��HMʾ�x���`?�AG�43��l����T����[�0K��Uү}�wsske��er�!��n�zT~�����&MB�p����}	�Y�.��`٤e������TyII��4�|���gɇ��dx�L�?�����e�I_u�P���3O�>ʭqi�|�s��'�~�Z�2���z'�,C5ndfV�;2���ۛrs�N�enػZ� �1��tim]��j��E���o$�$˴�[���Q�^=d_a�c��Z� �	�VEi�bKP������S�F�F�eځ������ƚUTTcs���.7`��u�v������'(((.���۾��d�_�w���$5�b>�}��gGr��F{���(2�0�ٛ�@[��_�^:\&�0��P�g>���iI��f���]	�ޠ)�jttt��t*�m0M�͙�S����F�mi�U*�4:Yr�hdb�(t.`!�&? $�<:���^f��___d��Y��t� ��;q����M�L 4��'۪���I@��b�f���60��X?����Dl8�$��L�&��uP.���@o�<x�Gl����l[���(������<w|fzz�7d.�ilh����už��R��Y���u�������ŗ�#��[���G�"����۠�X�(c�Ƃ���r�?���I�D��(���h �������������P�V�I0�SjS��jhf�r�/|QPP<�?C��f$� �D���0�*&���>))��H�ڝnۋk*�ќD7�s��K�M �j��N��$m͝�X �eo�t����R��d]������ǿ~�3��nf����{��h�9�4��.�ۤ�S��w%�/�����M���MB�[���u��񺴭����pA�� Gh3Cggg�
ZW|᷂.z���!��?EBJ�X�i�J���˄3�ݤ����m��-.���S�,"b_�;u��,,�
�/�����Q�X�"�W��qe�
���l�8�u0̑#[s�\ڷ˒::�k�M=
	ğt����r�.]��HGhYs>p5&��� <~�y��^�2fN����mi����3�k-X���������hi^P��(���Ԑ���M	A� ����n��ډZ�@*Z����#�`�WK�^0��̸��63r�s�6��kK3;!��Eu0������9d�x��T��l��û���C����hi�@l�ˈ4��L7���&$o����ɟ�����4 z��� yk���8������Q�D��
�j�����r�ᇯ��Ê��4��@�N��J�|����F�prr� �iYYY��]WN4���R���ԏ
R�b�f�?C�>"kd�r�O��Bz5R��A�*S�5�CrK��/mi����W��:��x	�'��ހ@�}`���#�����ؾ'h�Κ)��i߄Oni��;ԩ��r�t��3t�n�J��h^[&��T�y:��d�ӧO�'��d��b5�Q�~����yJc��o���إ̬,�dbC T�M�Ep��5Y��%��UT�a��?A��vnm�C>T��ߊe�ֆ�ñ��I�$Xmmn��(���J������J���Zi��~d��W�@��JB��޳s=��5<��N����� �S�Vd(����}��ɜ)��[`�K�4��b���ğ�3�Tf�d\G�<�� Q*�m�N��[�nQ��%������==�*`��h�BMM-<P�ܳvR�d�P�FƁ�7]�""X���KX��r��֖��v�����C=H��$���r>q�p~�,�J�?Ґ�V���.jho{��_he�y�ٴl|�|x<#Ҧ�5d2ϊ_L�@�;ƾ���"ߚ!�h��3���u��߂$"��tV�����@�a(Hϐ�_r�j*��
���Cp��V����ȳ�0p�9��q==��p�1�{_]�X�Ǜ�2�_n����+���l{��9�m�	�P:�oE����YɃ�_U |`�:L�̪֘7�����c$r>}�-���up��k�r ���c]5�D�>> QQQe���摏�w/nv&d��:#�a��;F@��O�^N,�]YZ���e�z��$y����ܱ}N_����M1d���[��A}��Y��@���V0K��H/7�d11�����������C�,�������̐u��$�eR����ʲ������4��m���ў���m�I@�:���:�@
2�P�LKK�Y�T�4I�Ίz�f����W�[O[08:\�5�'[����B�Н'�I0��v%�e�+�:��Ob�322��_�!t}����u��FU�ƻ�A���l0���/�I�^j��{ޡX��¨��.��b��֬_���Ɖ�S=�`�x�:���\w�����Z�+V�&~�b(�C�<E�U*�+�~��>"q�=;�gW��P�l���.<�/���If��ϐ�D�;e����ͷ�f�D��߹�F1��ˋ�=��G��1yl7�`i�Y�w׷������Α�?��~jBF�m���qc4�^��O�y.T�>�SW����h������F�o��Ta�P����oo�}%�~>&��z�7e&d2X+oYZZ��E�zF&l~f?c/F���_=��6���S�<�G��
bBCC3�p+�]C�r���=����@��7$G/��`�8*)�k��ڶu�d�\�!;D�% ,8���g�*� �g:g�'a�NhY�X�l\S���)�,=�P�[G�P�6�PSq��F�����"�QJt>�|�ZLO�A�}�p<`Okl��Μ1ϖo^�N��y6�S��ꭷ{R ��k��S��k��g��kE�M����s�Dmu������Qki�K���N��3nڏj*;S�	��q��ʺ�&O�e�}FhI��5�:�)vSY>Ǻ6=:�}c"-,�Y;(c��gi_H#�qP�[�/���J|4Wx�%��F����NQ�-9�L��-gާ���^ յ2�@iU��}%��M�;��8������;�P��D���D��V��o�JT�o�F>��?���^m�p��G<O��Hm	]�!�\Scۑ���|u��<k":�c�i�+�i�PI䃵����ᬂ�釟[w6�>s8��x3R���D�0Y��m�꧘X�OY�*Fe��D�A�0�dU��ɗ]�:$4�b��h��f![�����=�M;��=����/��Թ�˹|xy��Y=L�����$�[���^c!�<�$F~?kn�z���~s!�e>�q�����:s��p�y��'s㩛qSLS{��Rm�p7t��y�߿�9p/�&S�l͜�Tz��<e�>��09u�+K��_����~������T7m���h��-t(SW���}�:/�!�$���i���B�Ģ6s!Z��-�8��˗���9�n!D{�I��-��mڲ���;&��6ފL/''G\��ئ�x��������!��CPe��
�nd�e�����?z#HC�[񳻻&���-4"BS�:������b��2P��mc֚�Q�����(B$�>n�+}}�̣=oK���������k�"e�0��k��?g���$ւ�D�|rK5y4W{��_%�,�������3_B��8����@��@N��SF������Ҿϭ�!oZl�S�J��n�
f����A[@���6�.��\��g�����^z���o�E֧��#޿�C3�-��W�q43�.۶y+�p���{��#|�m��yA��������83C���{�i�5T�����䝣;g�n[��؀c�B��3�1��-�\�T@h����4�Uj�"O=��>�#�T�r�p��M���sn*�eJ���Ȃ@�BZI\>nf�f����4)6..먾�ܳ�q(�v�2Ҧ?v�T�w����}KT�
������n2�mn~�?���lz=��mEEŒ��,�>��p<�������!�	'�L�Yo0*yINV��64x.�G�f���X�+d7f)u}j7\��\Ӵ u��g�]*N��8�1z�o�k3R
�%����4�=��_��j��<�����yV�����~�[3�ڂBQ�}X�G��	:��fQ�Cb�Hn�C��P��UO��WQ�m:`�4Y���G�.Mr��������Q��O	�V�����e�㮵�*�V��@�F�)�0��縩��A?����Yn�)!�l`���/��c���buԡŵ����_�GƦ����օ6��n&�9���\58��w��Yo��&b`+���������4	Z6Z�����+���� �w(���Wj��\�u��N�������C����{������sԹj/[��:��@��C��t��#��*���pm��1�-�C\��0���쑉�?KF�L4Q�0����>�������4% "re"���d�?����MC�D�A���H�v�#?߃&��{��o;���)�?�fq/���>{���)?a�P�*����Ä13T�^q5@�Og���H1 �zt
���9��MD�A�'C�x�%�mҺ1��ϟ?@��1%�h]�zUbO��g] �A۽"	<{eL�Fs0;������AA>�O@��652�W =�����ɐ�6�o�E8Q����!�mlj�;v�D��M����=��h�<�s7|���͔�����J��=Z�nV��/�h���AO�fgէ���=�����_|��8*���v�xf��`[J�3J��������������������Q)mo�n2$y����qS^%}���@�_[uX�'^>#�j׶]XGٛZy�t�VbkW�]�;EC�Tr��ٹ�� ��P�&��d@;y�OG��f�	����bZ�.	
:�&~lSS~QN�Hek�t����^�
�DV˄� wo�����N���xy�l�lFU}�!t��Yq		���:�,��7 Q�u[�Zr����{����Wr��@vO�m�NF�g�2�5�<� �74��s;w<�@�gn��݃):�GRB���P�9�4��$ pݪ�Ot���M�Q�����Dw���x�K*[�K�O@��S���HG{�m!�K��Ši�?e�xP;O��O�\\��z^�(:L:3ohkk+t�p�b�1,4��Kνw��3������'�?{FFz�����3*�ުyDS{{{��q�<�H~Jc�W���wYXY�/��Q�0�1�z��
fڃ�qD����+����u�*|�jب)MQx�?΂�X���o~$��C�}ra�"Y�it��ׇIDޓ��ah̏�~��ݻ���Û�)L�,��Ϧ�{�l���'x� Y��G�PG�V�CCNJ4`����L~���6��K�T�C:������T���q���	�m�O\�qM|(�yћ��@��̐�N��j�����Ӵ����5�1��f���a���������W��Τ�¯J����a�dW�Ж�Wsp��N� �����+����j���#�L�-,,��P LXOo��o�E>$@�@s]����'�Ḟ�7�����Lt�<K���~��z�ݽt�����r��x��ϺEm����ً��XHZ��ɐj(u�>>F�|�)TV�4&ߟ?~� z����0p�'��۠�����x�f����O�Ő*�t*L����E��k_SP��>���VG^OO�:�����6��v��B�\ �2O�^N�6��*ܮ�gH�682�a�Yd߾}�0�	��ૌғ�M�ǂ����_�45{6.Q^���˷J
+�~���'&N4��ƺ�v�f$���eGGG�C��ʖ����������ѺY8r�����솆�
�k$�l=І��[�B�G����b�q���ܖ�S�N�x��,��~hu||<�_\��:n�ʅ���~M�u/��<�r�R�������乍^�'l.T ���㾺����Rj�Sk� ��t]>6xN穙����պ��<����E��$����	����7B-���ihO;���.�j�	j,'��� �'�hN|��'X�ߌ��������u2�79�k{�p�44�����T�PV; �HB�C��@ͼ))	��!����8�n� %0�8�>7���mj��1wU-�'x�E�X�
3�g!>>���$��L���]p�"/.Ϲj3��ѩ����`�s���bl���5h�K0� ��2�D�L�ی�z����s���)9�%��ڃ��$˵p/Q�,�p��vG�H~`+����>}r@'�t��E����
K�f�M��8�&��8�Q`ٯm�NHB৥�o|-!R� �*�Ȩ�vtT%�rd�ύ}����|��X�����C�̓�P��u����g܄�Ms� ��G^�I?PSS#��	=}y팖�V�F�$&u���G��SS0�@`��lįcO���֨ݺu+ r�l�z���{@�)����:z�����6��eeeZP%Rs[��FйKr�pz�����5�$Ry��QbRSyڛ�gwA����\�S�L����o:��3Pv?���P-w����hhh��d��3۵�����[W�0�V���c��QOlA�8�K��g��FILФ���M(�'��E��*�rrr�����]#c��W�5j,�K|3`�B��ε��>J����̮��k(ml��+�
�����s�p���[��V"��ΡW�
l�b���q���v��,L-C_N,|,u�=�`�\�|<<������z��{7��UUU�:�f.]�́�V����.��R|'tx��dv� 5e>����+=�72�W��S�jfk�������i��x"�.���r��TCC��9�bRf��~��Ĵ���$���>���\��\XX�y����63;[�% �ONzz:w�jFyx�O��G��������h[p�x'��$����Ycff�j�Ę}����q�um��_���N��{vv�G�ٹ(�^��-���c�����~�|������;���ⓓ{����`TB  ��.N��n��yu�;���H�v��qt��=��*��
:����f��C"�2 �h�Li�(7���WTQYd�'7R���BCB��R�v�׌�����F�����07�g��u�0;Q ��5��V2��	t�lm�-��Bb��Ĥ��ʓ�mR��D�X�3�X6��t�u*~*9��.i$��M��,?RUU� �9Hy��+�稨�hN��@/�$��Q��\�,M��#!���yʀ��&L�~�3��?L���{����S<�bU���ʣb`s;�6����W��B�;]P�xKQ�)	���c�kv����m8�}������A�9�V��e� 5�%Tk�8���?ߑ���F{�V�q4s�z]j��!�!T��_.�����a�0�bg�ڷ�2bQĴ�������7y�sҮ����VŏY&ȱ
�U��T��pX������T�]K@ۘa�.`���`L�)�g���'1�����^s.VsO�f�_C��g343k�S91���5_C�m������u�`��Uz�HV�����z�x��+�$��x��w���?�,�#�X���ؖ�JȠtbu�~IHo��F\;s-"�ݻ���Zw30�&�t�O�K��ڼ���(ݹ��?���ջ�@:�a����nkhP�[��	�y�l����=�؛�v���kd%zG$�j����D�9���G���>_��q�
Ŏ��{�HH����;��c�	.��=Y�"�\N�8m�g��WR�A�Ӻ�0S��g@$6���w�X׋�k�#ebb�����痍����>z�}�;m���#��'�YM]�l����Y9�eHcJ����J)+7���Մ���A5f<	B6nx�n��7��ξQ'��v�~���h!нnF5���=��l��B���'�W��i�L�,��Y�ʜ��,��w�
&5]V��Igv�MT�\S�� ���˝챡���S����N1�Ǹ�wEr?�tz��2>�|��By�Wq�]J��MDp�ܪ�����~�����ѥ��dF��U���ӗ> �q���B*��ګ�β�\�;�n��޴�X��L��vG_���?�o�;����v��~���|�\���M.��<���A�����������J��ϿG���4alU�׵��v�O���906�R�&+��Vа�[��6�I2��/��^���^BBV1���n�F���e�AOI��{���:י.:Bp����6��ù���'Ũ���<kg����Ϡ����O
�Az����&{:p���L�7�ZX��rm�3��hC��A���6�7a-y_-Z��\�%&��T��J�֫��~�5�˃�k!`(��$a^}��@��lœ�<]�ݿiΞ�s����-NWgH�?�>�_8.�� �4&�o�� ��������$ r�Z�ʤ�<a�=t�hZl�0���Q4-��M%�(P��EG	�>R�	�m$mggg���f]�t�Q�IO��H�*A�#З�J���:L��P��I�T����bbu��
d�s���٭[0����d�T���Wɮ��1���־/u��a�R�Z;��rd#V-��%��*��Dg=�ͺ�U��'ƕ��D(���R� �),��W��X�&ί��w���
�����Xk"��f�4&,d�A�"r�5��9�H����ݛ<��t 6��.�n�땯���_��'I��H�jq����N�]諨�DGF���M[�����D��Iqt枮e�̲�+%1!A-���kX!ꀸ�{�	¼T����|S��Y*RS]z����M�J���6�:s!fu����ѩ��/��9v�)�]8�t���L���e���7��$��M�FV'��i)T��`���ӅJv�K�V玩�)rt�KA>��a ��r�Z;z�hZ7�Tx2�|�W%��E}#N���2���p;�&EHrZz</��J+5-��u�.:J5걱1�{��w~Z�IWA�"�ozR�W�%�ݻcRRn_�p!S�����ꪪ*taS0��Y�ȣz�/S���̧��QT5�wT��'�E��y���=���mb#%&�7��6�����d����w��s�b�Z49n<��X����(� �łW�'j��
�~��3��mȏ7�cu�Q�, �q�%���q�&r�=�d!Qg�
��&?i٪���F�,%2���#ɚt��D_���[A��PhN��Z�l$�+'�tmҩx�}C��X��@y9��h�(��;P��厪�]T������_�'Ȓ�p���?�~o���$G90;;{�y\�רycYĩ������J�+:OMn�2~��Կ/�� #��F�A��A�ɀ�y ��W9���.$��ʨĖh�!�;���f��K��0T�Y�{�O�[�{��K+��X������gF�o�}���/�Hv�a�.\w}�_G�s�`�:���1%Z�����?�dh@&T���5��H����C�������K���6;C=�*QMu^[�9}������;������x%��'��Wsg�祟>��U=oimM6j���0�t	G#`Ҏ.��z�uC�@��t7�Ws���!�./��t��bl��~8���Z�m2\LL���8\|�qd����{.I��S���tHA��_��ט&������oJ;�P?�0�d���;��B�C���6���N�8��7�b���P����t��NB���B���kM���Ҁ�!���Ǹ�����{q��Qa����e��bH���1	��Gxq�.�=9��} �ސJ���ŉx�V0Pۅo�S
[j���=깾��lC|����/�4�焄���|'�~����@(��@,~�.�����ꄸ�C9&��^ܾ�i|��I����ymW�j7{�n��]��Ŭ;1�y*�����"�]�������|��"3Ur��AV �P/��'����=�m_	C�^��
����3�h�ݐ�=s0N���)ce�$���]Lss�c�𷭭�+�3u:�t��Udee)?�	��-��{ŕ�V�T��Օ yi��<r��5n�wEh@�����a������Y�K�q>��S���@��pLW%�&��Y�H!�,�`�1��1�e+1�z������0W�����ٝ�ͤ�s�ٯ��yK���#.��(xx�`��tp�rU}�]���z��� Ө�Ǿ�N�n����C保Bd�T�v�3r� �^�<�*e�3�3��ֿ�#]�>�O$��@�srK�"��޾8X�г���yE�3Ӱ)8�C���"�GNq~������hw����Gt�C�y��}LLhߔM�E�i�A�.���H�"`� �G�_>n�ϝasY�c��s��ە�0�w���W���Y��;�[��͟����s�*�Wi���Lp���t�4(���i#ło��=
��v|���3 rj�r����"'��g�oW���p0�+Rk]����	u,�
��D諆� d@𲽃X�o��o�c��΂n�Ѻ~���4�+���N�R"�eݎDy��;�9&X��r��C�F����\�'���rRT��}���-=�z��������:�.	�|w�e^#�|�ki�^�_�+��}Ļ}�����:�0�U��n>b��%��~�'��8`�z��q�R�mieu�~k��p��ȩدGԷj�/�VE�Q�����^��z$H����~������\�)�"�Py�]0+^�	�{@)ESö����ǎ�OK=�nD9���Vf��М���X��E����l���u?��Ǣ�ƿ
���|�j�fVTTD7��\(3?$�D�K��SY�LK��H�G�OaѣqC-is]�\���%�{A�݂
񧡩1c\�.ҳ���.ں�A��߫��p�1��F.Kq|����4�^&�<j��&%0��Dı��S��Ggs�����؈/̥���_�v�����;�]�LX܄�>S(SJVgִ�Ǖ���Є�s��m6�x�Z��3ӿ|12��I�gJ�%`hl�T���AnSb�\>�� �F�\�d���K�oP�WݪŊU�Kc0�֖�Բ��zً������v(�Y+&��?��N����L۵�/��0�ݙ�����ycF��O�vz?���hn#�����>==a�m���~AÆ��Jؕ�Q�8����֦�D��R^Q1��D3�ܞ9�ৼ�L���^��g����b(��_w3��4%��MKK;O�i�V��P�s����3KK�.\��2��x�w'�X�*��V%�qb�<=:������~{[��u�+:��)n4ջ��ː�k���B�+������*R�X��\�e[[qa%0�vCKd�/eH1��c�����H	�>cl<Dΰ�
Ω�僱.w��V�;9]� ���,ME°�C�6ﮏ��'QއTU?G埐�/�Ȝ��+\��X��w2����5{����hH`'g\�E���zg��R�ʕ����������+�q����{�`���U��Ѡ���F�k��ms<ވ��a�C�o"�.�l�Aq�����,x������w�ZU��ɣD�b���Kqo�e�Fw�9�A�m.���0�N�e��*tBG��!F�2���c)�0�?�K:Q"��ã��p�8\Z.�XN�h�S�(ݍ���V󠳫��\}����d�5���i�^j0�tk��O�S�ŭ3�a���p����TK��;���|ͱ�P�2�\�̊kpW���U0�Ĳ2n]K�c/p�ى�ۣ����m��z��I���O�ѓ�4eZ{��=��f��"ܱJ��lz��(O����Zև�j]�G��v�mmB\���5>�2X�Uo�D��`5�� '���Ғ������Bw��� ���z����IA��s,������TC��o6R����ʆ+:��<��mY���2I� J���fV8Ǌc�a���}F���;��f���3Hg�]V�mw�[�3첏|��\l�t���w��߿Wo�Ud�������k��?[���Ww��o���G��!��e�ZS*�.�͚��T��	M��u��Hu!k�%F��,!z<fw�Y/��C�0N��imW�b���U��YvLI�~W����ꭣ���?Pi�	A�k(%����;F:D����nQ�;����y��w����r��3s���s���Juuu���  emNXbr�x��ߔY�&j8Z��/lmm��7�����$CI�2�A�|��h��]ώ�kr�Ôp�0�V7��v����c���Q����v�2���`����u{��_E�K��Z���-�}
�7��\>�ÿљ�s�Y4��{� ����!�6ݾ��x�m�2���H@����5�7thAE�c������!�<0�x�4r�2+���/~�|	�W���Cyטx��3���r/���$	�������`���wA�����.b���PX_��n`�!۴S�B��Y���)x��T�]�>���K��⤧����2]���f}��Ye=��Mt[����<-- ����![K!&� ��r���0,���[����W ���.h��M�F��Ѷ���Ty�"X���ҟN��-�*����������a�������sc�-�>�.
�F��[QK@�Ƞ�hŽ��c�Q,r�mu��X�}}]�cî]��8-�8��N��~���i0���L<'y��,��7��RR',����"</��^�S�U��3��uVPT4b�kE+����}��R�۾���O���D����{�AH��~��b
�d4�8�@2�p�!V'::ziQY�x=|�7+�Q�χmP���+�������}��"4cc"d����Z>k��Ge�L���N�n����r����^�z�&��#�\w=�6��a�8O�yĴBES�7U����l�}�"�!��0�W�1�����1�;����P��\��Ґ��򭍗�0�A�U=&���a����Ͱ��/�&��_���ʽy���%��a����
�>U;�d�v�{`��/-P_5uu,e����L>6_������Aae�j��r@e-����~����d5Wn��sc �b���t�b�W�
�c1'�,�ڡEЊm��43\�C�*�[�u�=� hҚ�=���qm/^�W���C��4I�Y��m���n~���<�$ro_�DB@��|I�T[r)w��ۣ������"u�P�X�ӯ�N�g��V�'0���{� ��[\\���l���:��i�E�յ���d�����7��myz��QkK-l�K�*�!����X��6.:�e9����.�G@2z�4�W:��:���ro�c�KY�QQ�u ��0����]�l�?)��r��cȴhUR��#�Ʀ����e�6�\7"�Z>����GZ}a?��o�n��[x�B'ݔ���b�[&/��q&#:J፾��/+��5j����C�?܇LUkO�*W3c?��T!h�P%�7nZ�ry�(\j�(ǣO�)�&��z��{�������s*I���AI�͒&u����Pe�i�m��&�*����<���ɘn�<�$?�
8\|lx�H�n���'2�:~��\�|W����A}��亁�Z�j5[N%�_¤�%���4�����S]dV��� �v����R���KN�W
��R�-qZ�Cݡ�h�8g[�G?ܰ�/���7/�ӑ� P(�M��-7pB�!�u�?>1!G�7�OLL<���os�����}ԁJ:�">?#��x���>᠍y?:9�3�X{!����laz�+P U��7�v�G��l�3��:�Bw��z u�V������I�� )�����T��u1��� ���2}F���4E��Q���Q���~����"ޛX���9H��6� i�<s���%�� ���s���Kh�'Қ�r��J���8|y�ݵ�Q?J��4$��3IѪ����!�6/_C���*sp�O�N�'$$<�e������uH��g�"&(�sP��WW�n����}�	Y4��
�s�0���;e��"���t1�9:��`�0|�֗㇮�Ӈ���;<N�2���m��i{�9�lP�s�Q�3(X��0b�ߵ�]V���P�tE�B~8V���[qFe�5�ѺCb�φ�O
��Z����D����дWgff��Z���;�|�O��شB.�:��=���xm���k9+ʁ3�Ѫ!�T>w�z=�����9�3�lp_�-�A�c[�Pd���79O����W�@W�f���q��0��/=��O�Ѫ[\�۩��GM<�^��F���.Q�G;�b�rY)�����ٌ�㦙I�~�3��U&����=���2��>4�
�}������|�1::j�5�%��c~s�w~~^������ܦ&]������������H��8KFv�pv�i$���MW�M͊��4�O�Rk���x��y(���&������q�����E����֦a|����I��0j�(O<\��^w�t+���l"�7�ݮ=vr�N�22(�{�"_а�?K�񥢴���P�-��0=��ď3߸���Ӈߚ ��~_�;FF���XUh����m\�ɊMA�Y����K��Ǌ�������f��i��4�$�(ʼ/�
��A�W��3����gY����nϾ�mk�'ə�H*0���@������S�?ikc�ڵ"�����Ke�c����� �hr
��߿��P�L��sz���t�{
���Hr�ʈ�T��~�#0&e\��Y��]^��;;���7��~�������_P��/�.:������A�'K-�c�d���AJ�E�Co+�7�y�&!h7�g�1�^Ն',C�u�~��_	��_ܚ��mO���]u�s��sH�����/��s���&�G/�x�՗!��'��R��eNN|O��$6��G�>�����IQ��Y�J	Sӵ����G�`	m��딓�1偭�|��g�h%�Z��)C���X����q�{`��į�.����/cO��գ���!�m�$�۷X�L_ME��HZ�Nn3������M;��(B֟��{u�+,�S�-9��b�~\b1���z����m��� .\�U�<�M�&r��M�w�m�ױ��	��: G ���]�xƘ����l/�揷l�U�]�G�>AXN���Q��Ѐ;9(b�&��-�m�htB��r3B�S�'�A���\�w�v���?0pʪ[�7�a����&TAʨ�(�F�듲F�ҽz�����
�UU!l�N����}���}�kԈ4��7���nk�t����}_7�j�;6;_��*����XX�[Z|q�f�@@�#G�$=S�>a3~��0����L�~�#K�� 	���;��6i��M:7'E�:�n�"HJv�2U�ZV�� -i͞�o��G8_�`�?���? �os)���.��m�W�ڬYka.::��g~�~�U��ǽP�xD��J�����~!������[ɟ|2�7=����ﾼ?9m�C���}�$̼�.fXv���������ս-r�J'����3rl���M��K*ey��X�#)ejR��cS��ί_�q_��7'���$��i�'�3l>Z�1��$Y�ͯ��������G�Ao���|����M_'��K�ʖ��̦����Ș�7���h������Ûc?AZCOO�K��̀ ��%a��6vvz-f�q��F��y1B���"hhF�@^W� �t���#~VH�w������oIU}ܸ�B	&6�퇢���,��Ć*I��.�L9k���Ё�� 
�_L��\�9Z��\�^0��0�3{����B��M�	53���]�v�'����{J_�����
�3$l&�d�γ�^5���;ԩ=yXه1g���.i�����W#��&ߺR�f
��=�#�����S��hS��:(�c�z����k|���p�$F[�\�8��7L��Zg$$��T%�;���!2��(m��a���iA����o�zqk:*�I3RQ�f�I�0�>䳆�zY�Ȱ��Y�C�O��>�]?= �[�3�ܐ�(rl;����~���z�n�A�n+|���`b�� � ��?M2Y�_"�7Ra3��&�dr٥a�]g��h�[znJJJ����7MO��TJm.����h�$������e��@H{��[S��\�\�8���l�̂��wl:]��Uu�__�9CJ\�}����.�9�)�f�ŏ.&&E�Z���]��]��?*�0AK��+\z\���E��a�0n��1�����X�ǖ� )7��rC��������(�fLH�'�-w�M2��
�,Ѩ�.뻬�'چ'�y��Xz±��L/>7��3�&ȷi�5����yʗ�4!����c�!4��z/7�O�V9��K�����߾�%�����2پQYI�ׂ�g+�b�lr��/�#K��v"~��*$���i%�3%�*t:�[���Y�\�݆U���ָJ�BrD�\b=N#��b|�Iz'�"�τl�I}vXfIm Qo�pL
ҡ��@BBC9Z[oC�u?��7/Ê}�~��~��v^�?��&��ς%�;�F����a���/޴-\ʇX�5��a���ӧʚ�߷��u:���ݝ�'���� 8���W�^��Mq�δ�	�NnN.0X�WOYr����d#q0q��'6��|-d.����>�U����8<L�E1�[_wFǔLjv�Js�Kܳ�w�����pn����<��V���7褓��F,������wl�sk��3��9��VT�\�u���smoQ%��W�~�;�v���ٳ}��u���hyغ�S�#��Ȑ,�8����F�[��.�jK][ډ�"��@�7��-f�ah�/%�h���斖������}�/���f�d	].�[�27Gb�8̡��I-���}�$��X���e�H'�2e�NY�m����1t����^IP�th��$[��~E��etzqw��RӿaMڸۜKJG�W��[�u����T"$����<z�V�)z�Ns@(�*�0Fr����f���s<AB��PQ|rr�t��f���+@�>��[�3)ʢ`�S�C�d��fOb������{�}}}���4ٺzo�����7�2��%�޷_�ɹd�����$��h��E��g�o�Q�/���?�X��H���u@)O�<���^m##cs��"ܶ���^�������]�-��w�8f7d$S�%J V+?��)}�vwۺ��V�,�Z�����G�~���>H�DS����زކ8H+�Y�!�r\�j�3� {�3@8�Gh�(m���m(p����Zʬ��ȩ�l�*�J?��Nac-Z/Ts�D<��s�=����0�\�۬Ө��ӯ3*��.��09�z$�\<|��0X�Ar�����\���z��t������*q����j�j8��� �D��s;a��C��S���\�����%����e�5i�5����h��ܱ���<^������E��.%�#m*��wɘ�0���p�-����f4���]m���*�HSj��k�����H��}��ZQa�v��%Q����*�k���=��d�)-��8�|xshI"c]kL�R4�0Q5��i��2�Wn�w��W0%kƦ��܂����sA���;������'�v��[���|�-�X��N#LRSAH�l� ӥ�VX�����7���Mޘ(�J�˪I<�=}:�5R���<��2�\Ğ�zU��V�<;�ڛ��4� C��uZ~�K���:4<��Ca
o� ��[Ty�6{�^�S��}�/��.*UW/�����0���Sew��~�D����/_^@z�)�Q#"#��_B�%:Q��p����_�nw���O�?.��&hr?�f����Ar?qa*0�Ї�|U���=M�"��?�E`N�����>�)�c��I\i_��V��oy���B͙['��_�T�#�G�+xM��g?�<eG*ϣy�5����e?��6���_t�݆���}�z�$�m�'���8���c�~��
}��n��#��q�z��ȅ��;{ꬭЍ/��WK�&�����(f�Pjd��ݣ��jk�l�
`'Ҝ�����J1z�K��x36r�/9k%l�ƅ	{��!5�Q���M!!a�V�Q�щR���V���1���d�E������%���Bf��$͢��K����F��5��������_�h5�,��Z]]嗕�

sp~��1�\���tИ"�n�=�Y{�!P�����&�OZ'���a�}\|� �@B���L��W��.���Ϊq�?1���c7]���LS6��,e��fMU={�L e��ڂ'��)���[p��#�hg9�h��z�0�W��ZWjL���`�����q�@���g+��V��5 �b��� �:�U� =�W�\��Od���Ba�h�ToǂD�IO�n�^�d�����{҉?b;�&O�	�3tz�uXh4����o�*9ss����� ؔ�������d��B3�T�6��-,��ѥ,��P`�+++_y��x����g�܈	[j�:>�I�}���)��������87'/��`ӭ���j Cǭy�z�EJ���2&,�"''>F�E�����}��m��R-���w��ӈA����ܕ
l����l�Fۖ�d�?�|�)C�_A�����?� v��ߢ�9Y
�����R�:���~�n۾Xl����gZ!՛��������e?Il/���i�����=
3�?}7���X�!F��b�ѥZ$4��Rk�OD=$�vи��U�}g��~����j��'���5B����V�b��h!]���򅅅2����R0�:�������F�J�nάp�y�@�7��̉���G���L];��/~�EײEu"Ve9�@C�!#'�3�E	�C�Z)A�d�����8���Mq�d�q�c&ܚ�#���a�����>�0�� |�x��4�o��a�A0`�eD������u�
�܌>.�ԉi~_o�����v�AL,	�'4��F�[���l�
Lj�X6E.�T�@h���� $
��n9��3����(���#Xy��I^(��,��������3�E��d����;6~�K�k��P&�����p�[� �J��m	�/E��NOk�n����
�c0S�i�m=�b(��!������t~ʶ.���eo�)��sj$���R�p���e}O��Q�����M?P%�ՎK����e�4lrx���N{ڀf��)����#�l���fY!���&���T$��X(��Jb���R�(F���yf��x�b?�غzZ'����F=d�=pi,}���@j^C�L})S,� ��5���bhG'<�u��Q��#��п������~R�-]ː�{�:��F��^��'C�B������ͦ�-J���y�,����&�6�D�����?�jc�΃�.�F�B�҂���^g�v��S
:��F���3Ј���"t�55�띌��<e@醆Ry廫�����f
j�Ʀҭ���-�T�{����#��WؠSjDDDeHHH꿡L���뻱�T����5f���-"w!��W�I@�J4`��O��Q=c�%D�k���WV��k�Bb�(����˃��=E�8�K
�f���
�S�q��-I*��l_����ȹ�t�![����q�~�P\_na\�Cqe
ԍ����! :�_?]M�ȭ?� ��n���?	D2w����l��,m���]JP���i]��2lC�
V�V�g���n}jr��]����"oh����Z�j�`�h"b�����f��Y��^a��i���͛7_E<�a��-�:�Կ���҅�x�u߶���-�������i۹DsWT���{Ci*���~3��U>x��" �2A�������V���7�R�.H��O�P�@�akx�F������ϼ/6¢��(�0�9�>�hx�?��ۃ��1絜t�����g>��_�ꗿ�?��!����@��i4���d|���lu��rRd�Y�uG�u�M�8À�ak���^Ӕ���_����]��M�;��p�A#PXj��xxZa#I���<�.������Ic��w��rr�i�G�v#|9�̜v*ފm5��L�*�׏�{f/�J !|����|�	��-�����>u��緉�22&���*E��%X^-����'�=�Ė�4��e����}�IIIi{����k�f>56BF����m����Af��kl����U��O���4����?�y���cIe%�\�ch��s`b���X�>����;�u�t<S��yg�TX�*e�-����1�(�Q�z�k5��l~ҲEQ�j}�,��GR��S���Rv���J�W{����J������Q�S}�S��쀈*��-[�x.%�Q �v ��;���/%s�����8�@[���:�M����"�Y��6�Mp�"^IG�V����k�n�'���t.�����%F���42P��KH<�M���`�$H�
l�����>��ҳ�H�qf�+#��Ֆ����@�:�����"���Pa> ��)�h44�\b��^qp�ZYկ��/HflV�R������`�#l���1@Q�ۜ���7c����L���9�&a��\���^�w���g��L{iQ�K��A]�E#��3ϼy��U�y�v���<=��:s�Qr�(
�6Zä�.�O�Z >V5̊������ ��}f��N�♏�"���k�)'���\��lH�R�!-ok��@t�����D�ݢ���D����eC�j,�<h
�)L���5\y)�Ho���b�\/	���Þ�e`c�
D�!J_qc��洣3�oA"c���@UZZڗ�����rI��Q��Ԛ�K���dx<CG��Ɵ����������}�b�� ����OKG�v^�7�ncgםĦ;<�GN�2���W@�z[�y�|:+[MZ���36�h��~�E�=rWE��c׶0�dS�NI7���qkrb�)~�BS���w���ޤ���0ӎi>�B��Q���0��1�;ie���2��S��Ӽ@�A�,F�Hz�ΠU���$5���gЌ�($&u�����^x���0�kNi�8�4%�05���s�/��1�����%��ߘ�9RzȖ��r��wf�dN`���A�$ � $����c����w�L�l����_�c��ǟ���ή�@麰/����z#���-:::�rYjF4�%c#f׻�dg?�B����&��J��)p ۰�:;T#�o�v5I�Z��hO܀���������'T���c[&������Is{����g���4�ǘ�7[]��EP����uj�|�E��K�}���U�3_����͠y$�Y(J&8<G�smpQ$8~��">Q�v�D�t(�g��11b�����'��G��� 1x]\�}����A�N�Y�fx8�`�Q
��������UG��tk�sh��P���L���I>zq������H�9�8#��: �b n�=��*u��ߣ��Y_2|���H�p�v ��WG� �Q �����_�i���B4�$��mfwoo[_V�#��Wu�B2�!=���S��Q��j��a�#���9\G�wYfH�����]������/�+��%��Z6Q'���S*l���I���h�V�[(�˻W��[H�H�_�ی��QkSyy9y(���"�]�Ӄ֯��ՑϞ�K�}W�&u/qQtvsg�분)�r ���F
�/@��9�P�&��L�Ǟ��`�[�s8@.۵�� y�tdJ��<e͊W4���:��-@���l����r��lM��q��]�ީ����� ~�.��b?c�յ���rJh:$	��'��y:�&"B���,"L�M�0��=��=�gl#^�(uv��XSQ�����X�s|��S[�	wo4���c��X/�*؇2Zbw��9�f�2B5���[�/E�}�8e���+���������}������E:���f���4��.��/Q[�4֭�����C�9E�����K�ab�2H#=H-⇨B�h ��	6�g��1V�V�['\@*4L]ӑ���r�7�j�\ՀT�NGj�O��&@���k����i�'?�Z���B�{��=e�|��YV�[�	П�`SF�GBqoò��i�jk/��*�����@��礤��zzzԉ�/!����j"�uo��#kO�����
������911�X\R���;{Dvи[�����2''��xa��.��EW������7�hx3%�����!x@(�r�j@���j��J��ZT]FG�Fi�t���/w�b�i~��O*�����Jw�=�hG{����Y�Ͻ�u/��u_	���"�L��ފ��oz���J����O�����:�<��{x����7�Sō�-���&
�Z�>���3d!.�\�&�5̯`���o�lS�6�E��0�PI�v/Id�D��4�cϗEId����u��sf�m�*&J�Z$�oP��k�|{NFv���'������ zn!���"vc��GK��,�s.`Lp�V��g��Mp'�hxy�ⷶ�� �яFH@�L��
3��H�=�� 7���e��dL��o-H���K�DIT�=k$h�h�L�������I�ys1J i�{��f�������8�������L�`d`iMxԗ�+-�����1���	�`ʴ8���.�T� -꯰r��Y�ܻ,4QN�_���=p"l�������z��8�E8�Z�,
�r~i���I�'�����;���ˁO��*;j�eї�^Z8���	���}�-�L�<�D����a#�f`oE�;�������GDȫ%p"���f�؛A�c��X���3����� Ӆ����	�AJ���h������"��ww߾|��9b<k���ߛ�� $\��2�5��I�T�&4�)��׸��/�ß��1�d�ќ���?3�n�fN��gU�<����_}A�*��y�3�<�	k۸�׋�첈���{�v�b��џ�Fw�"�EY[l20��t��.�Ms���N3���$���Գ���Y�/1U�1 }1�gl=	�汩�s_�EjKEF��H_�p].�k��_��/��VC��#9�G����?wbH���.G&���"[MD^_?=��p�+((hj�Ϸ.��Pr�P>��sP��@4\#�X�+(�fd`�v�@z��qfgfFh��w�&H��v����]���?sc���`���������NYi���*�J-Vx-���H�k�NF�]��E㈊�*L>u'/|ӟ����'�4Y�z��n�4ޚ$���I�����3偀�}Gʰ}.*  P��� �����+���p���|H<%Q���d��Ha5��"�s�C�F�fX�	��-ݓ�^�#*��=���m�jA{B���a���������MC�_mD��F�Ksma4$�k�Rnd���A�Ń%p�d���F�Gw�����q�Eq�?�_�Eu����hZ/F��W{��-*e׋=m33��q͛:Iz �츸�@[t)�"d�&)ݚ�=O���-�X�8���<���Z�F�MIM�0�����B��:k�l��'{��82�,�%��Ñ��Ri7���Ņ��+$��גr��ψ�/�'2>�/����VDQ�^���*b���
r�q|�6��![m� t�dhr�:��h���XKǏ ���B*��f� Δ:;<�͝�N�`
9�,�O�� ���N�?`��2zC��㊬Y�~�QȻ廙;}�?�$� .z�@,	��-��u䝆��$�w����"�i#9�Ej��888�J����8�-՟>=137w�g���
q?���1N�ߧv#www��Y�.[�V1��Bᇩ�$�o�������Y�����8]kO����P�[ʇ�Y�C\Pk�w��+�p�<�M��)��X�B�hv2M�l-m�7
�m���nnM4�9���X����^vC�v��o�VG��-�2=�:��	���K�_Ҿ$>�@*­��ÉY��ds�J{z�����5Е��v
(�f1r���?�<t;n���2Z�	���a��c�S��H��9*�8��_�v'�@���o1h+jh��� �ypL�PB���~�J~w���-2���D�s�k���>}j|wu��_�|QŌ���B��zY*w�=��S���Ժ�41x��� ��\��S򯮫��,
[2r_G؛�"P�#�m=�|�=�r �p��9Ą0�� ?:��5�'������m��cf���|�Ȟ٧���bGF��{K�
t'\���M$���23��2��H����2-4��(�9|�����|�F	`1���M���˼��~Wj[�W��k(A�f��f?[-!�a�bc�F�壸��?M��&�wO�+��\\.N�9��xT��_i�-���[��B����'8*LNZ�(� fӡı���OΞ !����
q������n�22��B��;�c��|��#��m��L�� �jj29��jjc�Ilk�3SF�F�����.QNd�\$����6<?`*l>�O&N�|͔`�+K����YH��p_�ݜ��ZddW1�M���$��~�猅��)[��y�����M�\�@1��� �: �9�O�wǓ�dCqM�A�h<nV�x� �x~����y��~e$�_�Ǔ�������ϼA��~�����]kl]�+ W9+��=���+���者��9�Q��i�,��h�w��ʾ<�����E¹&iu�������*ƛ�]ԧ�lV�rq*��KZ��ו��$��]�w�����y@ˆ]E�b��9mӬol��찺�
����A��n|jj�����F1�������)|�2��K;+��(��̄�5���O���%EhA�����s��l����;Y�+����lM��Ͷ�n�>fJ����|>ˁ|I2e����ݙ����3��?K��|߽����>[�O.o�k׎"�W�B��F'���0<9�*��)}����3�x�����-��i�'f�&1�sχFM[��������:��A���n��qx�)}�K�{�6���,�KE>����bps�kG�I���weҾy�?���($D���*�Xb����Y�?��Юc� �>�
�0D��GtJ.V���o��輷`��-�gA
�,�\7��ۀ2p�Q-���r�gd�����X�	��	RDs�j9����VY�%�9be����U<�}e}IrE���d��Ɛ�>�h*����:�/vB�z�����#�N�o���[Pr���OѳI��8RS�g����~{����A���G��G*/q��ُ�%�V ��=>�$w��8���_���\2�cO��G�:�q�Z��;�r�8�C+�����T^@��	�s�l�]I,����-R����_}���ܛ0�=9J��[��y��w)�N�f��L���3�M�=��F�r��d���8}����o+��Կ�i�M�Hb��M�c{���c .p������YYY��q~(�UZ�+��u��09<�*����϶�daS���CBB��������C�)�����.�����e���dQ^�_�����"  �g��m\D+��_�=���f��X���a��=��
/�,$����5��5��^�����^���ش�z�"����C	���2�Zj���7%�S�њ5x�BQ�vW,~Z쐍F)Y�՘���t��S!��d�{����]���e\Y�����D�B_n�����۠���+�]���U7�l�?U��%�{G12a7�������R�V��ϑ`���L�f�:�u1��&��o�94n3 ��FB�ѱC�P;�x�NSRRj�)��᧓fm���\gĳ�C��;�;99��{�J�ݞ��ߤ7���3[m�t�ď�?M��ШI8�V���uYY98�s����w�e��<��h��[�$�T�⭳��]yxxEz�/�ӧO�63s)c�R22(�-<T�{��^�Ō-#�ft-[�T�*L��ӂ��>環%�0�=�!�~]�~g�c�f���i�ܣbo��Hؕ���aiۛ��K�F~ k����G4ʲY-K�Rgvz�6�8��yN��	�+)us�͝�ö[�Ei�A_��>�Дh�q�1��r��[�S?wƩ(�.t�� �����]�^�8�'e���Č"j�I�uWLrD|�PÏ�D���$ �&8��B���৯~����oVI�K�j&ͱB��Ds7)�R� ~̸��ߟ"B¨��S�	�mXcB{{���$ߙ����<Z�t�1|�A���#��|,c�X�@9����od׆�H!x�r�.o���8W�[��J�	�> ��Ru�P+ޔE��R����u���m�`��h"B��-��R��� �%%k�D���&�Q�!j�3�����v�T���Pճ��l�$Ѽ�ZHL�h������.郾:�r.?��.�G��tw6��t"2_�B	��ow���ۜ�W~=�,�h��+���M�H������ĥ����`я�����p���i"���o�mo=���-�-�p�_�D�5j6�D5��f�})�,�} �Z��ߪԃ8�ی���2z�Ɵ����,Z@Ԫ���ҡ��Cn�tTb����8�G�H4~~~�@��.ќ�����8ۭ��Q�ۂhDdd�㒘 Es�aЎY���in��H��' ����4�P'0�!��Ws9��U�^q"A�����a�Â���"�B�U)Pg&@��D�W/|�(OX�Z@�ά�U&M�@Q�dR9o���K�8$eo��� �}��YK'���aP��U}�b�'y����L6������;!�v1�ݠC��t�^�R^����չ�JQi�g�:��=�'}�п��Pn�nB⧷����'���P����M��ʝ��Fy"g�De�9t��>�,� �I?��_��-���c�h�{�����-ܡ9A�kA�����l�E�U���Av�v(����� kp�/3?�A�`iaOѓ�����"�ǄK�d�"��&H���3��eϯ�+�U.�>�"�B�ܵ�t�J�.W�����C�b�WO���I�'�%��E;*Q2�?4�>�D눋�>�F���ES�G���H��*Ƀ�F���4�~&�(�.���;]�Hmǟ
�����,@�Ӹ>�Y�৻(9�.==�s��7�-%꽮%"�p"��ny��쏉��%��o�=�X�@�d�� �t�7ՠ�&�E�Tid���x��N�;dS�|;D)��8��9nf_%�'���7<�!:�/ �fp���2�0_�B/$�W�Y���مσz<�FK�'�B5�`�1�~�"Q �)�$a�8��Z��g��':%�0�X��;���+(H�`��F}�X����롗�����!z.<����Fp�,��w����jk��joA��za$6�^O��g�^�����G����ԦHhC�t�Q�'Y#���(.Zچ
>�/5Gﴣ��m�O��-6�q��W�E%�S�!�.s��Z(���N��?m��B�w��ڋ��%�j���/y%y��BTgH��ڶv���K�_�r�I����l5%�l��U��s���Jn��z�������6������{���#�ÿ�A>=C(,,TQSQʇ?��2�5�0�<Xt��^*�y�6�'�jE{��H������Y���\��T<�-�,c��zG�p����<�,D�x���ӎ��gu�R.���ٺ�$a����+��,�[�>H�,��<ӹ�`+�o�8�`(�	=Z�������4w�X��Z���B�ʨ��9u*���R�τ��4��<��5]KQ\������<�rQ����)؛������?�רp3.�Ӿk��=j6��t��j]U財��;�%l�u�t�w)�M�i��RS4/���$ɟ���X̶�Ø�J�$��O_�/�dA������T^�	���|�+\�����c9Bv?y�9��,�;�}�2-z���YxZ666 څ��~���r~m�ߒ��@��1�,S�#"�Y67~d�Ж���'�ߧ�:���0�L�d\�����iӖ�Z�ӹvtq����2�E������-��Ԥ�h�|Z �a'�3����Y�#+����*ֆg���B�G���*ݼ�,_Ms���u���n�5w�w}�tm|�����_D�kz�4\4=����JZ���`�_���C��$����$�P싃���K�����ފ�W��R�_#��z��nymln҉�REJ�Y[0cj_А���)���d0( 9������n%:H�o�~���3�>��x�륟���F3-��Ĵh�t�����/DXhI�29���l׾�cd &<�̱�3����P��W�Yﷰ�Ÿ��j�myu�Yr��Z\.��ĺ�Z~Uf%��D�T�����]o�����T�#}�����vH�|	���:u=��H��&�q��*���M�1�'tst���['�"<����я����x�]����qo���m4��`~��Zy����L�;�>����%�`�IPj�9n,N�ml��D:<�c��,��ڨ�>6�լ����y� *g� �,NQ�/���*Q���@m��R�N�M�8;J���m>��0}�W�3���!2nn������XT�F����sE���v0b�p�R�>���Κ�x(}�X���7�w��2��u��;��A鲰z;,F��F����j> n����%���o���}��N^��F��P�5��<]~{VG���kjF@i�1�ٍ?�bK��2���/*���A���$��@��	��Ѥ2J�?��#+޻����B�#s����JF{�<[�����]Z�p��qR�p�Y�p�3�dL'�G���^�m���7G��T2d*D8�"�~H���X��Mlֳ����_O��|�]s�ͨ]��V4������	�+�*Yn�!�q��`s�ѯ���h��ӭާTR��s*��>K	�k����p{y��?]��؟����|�a�/�@�uvJh�hv����p��J�ptZ��537?Fbǭ�q�bR�A����y�oT�ޙ &1�}�`?��M��W'��G:�ͬ��Ȉ6;��p#,"H��:{��O����Q-���<��!����8�8��^�ϻ��\��1�����<���V24V�bW�=^@���/9u���_	
�15:D^�,I�q�V0����ꨨ���AQ)I	�����T���DABZ�[@D$��n��x������t�q������8����,���VՓ�%>?#j���f�wW���gz�?���ܒ�Q�%)S����I4p���g���Y�8)���z��M�5�*��[1����t��ӕ<�qG����ɡ��Ɔ�����<ڛ7w#�Eԕ��A���B�8����N(�*��z����~��R�Yn6H����:��Ɗ�b�'�	fo@`���3�C�X�'ƀ�d�r�c��09{
���m�Ņ���g�L"5���4��F��\J������LcH�RD��<Jz��Y���+���a�Q�>Ɍ�s�v .��]F2�䔥���=�9�MLđn��[�W�Y��u�/IZ��7����ܝ)�$���g����V�q�C�w^�Ȕ����`ëB����&��)n�3A[�;a%qڈRΆ�����_R�3��ӏii}dc"�Ԓ����ev�bC��@�)(Ȗ���$���P<����M���0k�j_K(w���2�8�G O;�O��Ut8��U�|-b(���������]_��~s�����dm� �u�3�);���`�n��~����`����##GMMa����&�fP6ٴ�z���4>�C�6��o�q��Ȼ񒯗q,�@��Ri�q��"�s'�����l0d!��!沅��*;�T�ę�t�t��Zf��[p�3���P������b�xxw�%��7������e��@g�|=c府�@?�N�������}��*;�v*-5��Y�o�.�#Ra)���q�����у~mzb��|�8T�{����#��:)	��6{i�ƀ7� �#���(Bʱ[Uuik�3%ẍ́���c�)�q?��p�0�c-�a���!�3����g��k�P8C�B���eC��-���RE�58�����q��ʓ��c���'��(
>�̝A\"���@.��^�4bm͔6��nԎ-<��n�&�䟺��A�"�G/���.ICq=)ᙢЧT�M\;}E��x��+ؠ&L�|}u>�n���#���v<V*D�N	6_��?�i	K���"�1����5���J���'K~T]!�׾���[}�ر~yz>���8 ��8a��V+M���;Wơ�`�U*)�ZJ@v9�K���E/��(F����q��߷"[��/k�̲U<��k|`��س58ʕ���+o��>��\�@G�$��f�;^ցR���_r�}W�*�Q�K%��v�Fww�}<<?_X�h����.���T�I��3s�(Kt|dm��a=u�Q���x������L|����"�k3�&b���U�F󡷣l��î�2������",���3��ln^����K�/�Φ�,C
�`?8kwՉ����~�g�̽�Q"�^��%<&�d��u3-�L�h*���<��U��o�@���i�r�%���:� �^�����4���9�f5!�L�|Q��l�-�O�Zr�y]{+s�ߠ5��"Lj��a=I��<<O��/��T�� ���D"�65��JK;��?&$�I��y�R1n��������J쩣z�G����m1��r�I$0L����Y���̺�=���+��d$�A |у���-��*""�l?��`[��X0d��j?(iw^[yn'P����)u�_v��UX��u�����6O	�5�]�����������	��Esu����^q�2�'3O��+A~�*lGԳh�9%���4�?��R�$����FJ�#�a�>ߔ�U��L
��#/*�~�pn�3I|,,�2�--�G��9_�ES���ݷ)j��Ds���gTÍ�[��v��x��:���T�@�k6R�Xϣ�Q��%&����]�hʲ7�(�!N!���N�z��=�������x:!����v�Q��C֝m�<���|Th��l�wkw����;����n��G SA�]��}^�.Ш����-L�����A�0��!�ى��S�z�oEruT��;g��װ)�?��)f9Y}��e�C�)A��qbbb�ϵ7�*�N�Q�����������$�ת��k�H%]�F�j��&/Skk�7����X��PX��l�0(Ƹ��^���^�W��p�i)�ܢǖ˭;�2�&�vߘ2�K���9~�8h���JF؍�>N`gWV��['���6M p.ۨ�
�ZT�$l���q�멉dm�[�!5��s�vME��M���b��ɡ[�Tp������X�Wҹ,���,�i�;3���T�C����e�G�=���8~���HL�hA~~�H�6���_��Se���v;0^;r1SD�o�����f���K�n������NX��!,��UN��O�^{k��>�uT'��c��y��r�^d��w��;f/"�B�f�l)*�g��΂��[~�z��[_��Q�,F]��PԷ������5'=��e�N�M���y7�j�����p$zq��R�,�߲�iXG���	� ���/�ҡ�"�H��?(����Mt��*��/_:��߯U����A.�����Ee�g_a777	yyq'��5b���(���J��?V^r�u&���[7��m��o���Ӡ���`�{���~;�w��
S�r��ul�S�s����7+�÷�a�xt�t�n�(5��f�vx��.�{; ���*ϣ=G�}�~�#���&1-o�����o����9��x7���鷯e�p�_LceKQ��lw(�x/�Y�oߖ���`��1����5�z8�-6�Mߋ�$
��Xd�P��9u��hck8e-��n���ь��K#�w���G�ʧo�'h��{��%%�t�����Q`���*E���F�
f�Hrr@U�G�;��� _�b��֖�@+b�����p�>8Vi�+%%5���r�%��ʦmV��5e-�a�#a�p�lX/	%�ZT�������ie8m���ۼ5l��ƅ�d�[������o��	�ʘ��-���BTz�0���M_��f����if"]���h$p���oK]7y��*^D��ś�xE�E��x0���:����5��O�:"6>��6����߉,!	�n�D���`?6v�6�m,P�����Q^�'KS�����ЇJ���l���������[X��b�~�Z��E�D���y�����B]��m��9��/X�B��[���l����H���̢�
V�n{��R�R��̒j�1aI*1�<�d���ckw� �I�j�c"^�/�k����_JJ�ux���~�҈If��O���J�A� &�O9�<J2&�`�i�ܸ���-ѣ��U}r�w����Ty��<m��y-���]�gP&@6�>P'��劎�x2�^���C2���/��6M�ڏ��"��Ԁ�:f�%��p'�Z�@�Q�>#�u��#�Q����~!�i_��i�:C��E��51t3�2�o�/j�f�lx'�e�N�Y˒�}����i{���CSS�	K�|(O�3�w��*�
y�N��OM��k�~���z��a�ٓdJ+@_�0�ى =T�Z����tGd���ng#�LrVgA�����Wl��B�T�]�^;;s@]�=Q~�X~r��rX��I�zM��-��� (�uԄn�z�a����ù�MW�p��e'
w���ҽ)}LG'@���.�
 �2��\�=;h���)�U���?�z��"����i-)n<�=V5�%�a���ܐ?�'q{U>bVvh�H{�k���"�;�����W3���B"��t~��G���slg��{P��N�#  ���i�KLr#��䠤����S�۞�����P"�KbNNN`�+=I܎4���Ӿx���2�U9(��QPP�Q����`��R�5��i��\(yU��a����ߋ�w�6�����B���\������}~.��e�p�-�58x"&[1R�W��RPI���Ly�v�!2�nj�}�l�5F�07=J#T�\.Uכ��R��*���%=$���sM���iO8s>�Ѵ��������S#���F�6w���{��q�6(��@�X���k4MMM�*��ܖ����L

��"�����&�~>�
�1n�W�-s?2&%�͙�":b��_�r�L?�I}�b�>���~Q�3�v``���F�E��t&Y8��1^��	��D�!���g+2×�U�n]]M��j�A%X<�v��^{xEw��&>��5=��1��BLd��Y�O�[��@I��ӈ �C���fI��?~�n3��_5`��M����d�^#���vF$����!'V�[���쌸Zz���X&&qKw,CTJJ�e��T�===\j�Z�8-�B�DD����p5"����;	_�@�z�0z�~�`�A��)[X��?��$����^�bD��QѦ��X�\��J�TQ2[e��F滗�G�ܳ}Z����g�i6r{c;���\UG^�L�0:��IT��l��o� ���}�2������>S+�.ʲwE�$�!\@0o0����6/�v���)�'�c6�O�z��17��餅��L�ފm�%d����CEš�{��h�*��f����1]v"g��K��j�$r���/��e��"
z]6��&i��JCi}A�T�Z� �u�D�ah�}���|G1������%�vK�iߠr����cF��00r�8���M�Y�?_'*#�2_K�jG���S��&��q��[�DC�m6�U1��/�����JYo��w<���3� ��������J����u�v�C6�.�(k�6f�"����|�C�!g���ǰ��O8��W���3�qc$a�Q�<q�����0�N#�o�㙮��|6Q�}�k�b���f��Q�ר%ϻ�:�>�j(4`�[Xx=+>u�WH��d-Ȗ����K��������o��6P�?��PUR��:Hs?_�U��*�����=}p���u?$��e5�^C��~ ]�^D3�nDCt�ӱ�H�@���zY�J�o��0�����}���I�!�Ϭ�q�Zܦ
T�)���&5;֤�+������z�Nr����G擔�
�(=$l����7���VWQ!����ٲ)8��M����a\5�AUfV�co&�.-P��lQ�h�������X��w�,���������*�E���j-��7�V
iZZ����rY����6���ݻ��xߙϡF��E\x�Ul��D�`*�I���SrV���YVb��T�G=d���%��:��xÖ�F$�0���1mZ�u�v�8S�	�-[��c���ԝ�\��SЍ���U���J�X��|�DG��bS�k�u����P�\dǬ޳t}@Vg=f�7�Q�7�Ф���q�T���tzAȵ��g�Jh.�)Q��y?�"*ؓ?����n)�L��%%{���3�뵟?����Xm3˔��Q��C�1�f��N��o'�iboik�%����'�an>9s����n稈\��w<Y"���F��	!��l.��Wg�C(�򜒅ٶuK�:Jbh'�X�3�ޅ�$�+?Ϳ+64�͜8�G+U����x���i������Y7��EP*s9եz��M���l쪚n�\�o%��=�@Oy���Ҧ��EC'C�����RQ��xLRL�e�ӋL�!s0yD��*�\�\���-Ӷr�`�����u�aH���,ӧ��^U[��GUU#�lB��=|M6"U/��j��'�H~E���t�����[Io����� ��3e+(*zѽ}�����j���OUuu{Љ_g��{ނ'~�sIS��J�L������DfXEQ&v�-mA7Q�Y7�@Lگ���}��ݟ��'�e*�m"�� ��o�̊
���^G����_����7�����_T#и���k���kQ(��i��w�z:��$����]���hq�j�j~�C�(^N�!�7Í��vx�q`!��/��T��[%�_?T�����rP��r��q�E�l)`�ƍ�5)),���ЗA�)�o֫w�RRV��!w�r�NX�C9VP[AA���jltt4��oB�T^��2;�Ah��?����}��I�N�]#(KS�����X�/C�z�źd�e��P)��#�]��{V�_�`nƣ��u↤�ݙ�����u9���N^�wihZ}�����NӹreP��k�A�BE2�{e9��DkfB�7=�/�Ӿ
j(e�|/���l�v���2ő��KT8q���gS]kX�>3�����g�X9L#�/+��C_�\e�5��!��EH9WNUH�ω[AZ:���[�nu5���'�7t�%�_�]]]D�Բ�Y�J�.y������ T���XAg�����ݜW�U�i�coG�H67!_��v»?J�Q���hM�e~I������{�˂"��>�~�=g�H��j��Fas����1`a��,N�
T�7�P!	}3��]���b&1�Y���sם���]�Ɏ����8�����JCNIzr��ȕ��j_9Wf����������x��8#�C��tԮ�d��ǰo��Ǚ���2��$4�����
k�j�Ԣ���Y8%QD��I!<###s�e{.�[.��ӡ/gUQS����}y�A&дӺeo7����:1�5<2�����I���O�Jw
��3�[�Z�,M�)��=6ֶ]V!C���+��?��Ӟ[J�n�G>�gS�=6e�^w�=��͑��Gi!C�6�s�G��W4�6�J3��*�tF���d-F&}�����;%�U�J}�3XTiS��a@8y5V3<�cH�H��Uy����ƽz��j]#-���6�u2�FƂB���ק�j��چ9��d��jj�X���ӟ)~r����T�xO����˫��S���^`��M����h��r9g=?a����b����e���cP[㽮��~��$|���1��Hv�%LO?��}��A0T�Y��ьs�5�*y#�'�,����$�`��#�(}���gSV�z�ޙ��Y�n�H����on��7b�Tj��}��S���dy�t��9�g��`?m
�+�+�@u�S20��˩�Iސ�jaYޣZ�|�})ǃd}�B^gD����j��}4 č���1
�/Jq�;���o�^,��ri�'�
 b7�	�I���{�Y\,�W�~��=sSS0�wqM`0�-�+=vu��]0d<�<-Z>�wQ��.9�����y�=^��vC�0�zp�/�F�iφ>�V&s5���`m��V#��Qj��A����3��M�g��M8��_�Ṡ�9�PO���~��-�Ƹp1ʉ��ҍ$٧ �z�ۼA����7 ]]֨�i�?����SW���r=�Gn����<�d\�ڊ�1=;��c��r"������=V.lffFOO����u����yͤ	�u@�v�����R�Ƿo��9��x�i�\;:&5uFݙ��oo���! ���Gy�x(��Aj�`\r�g�bK�R�X%;��B�����=zgd��W��I� ����If�^��&����H�fw�xs��d�s�>8�����HOe>�^:)%!����0���l���IC�B�Þ�u�94*ʫɣ�ӌG�k�Z��i ,2"�o��&e���j�sw���ui�SM�9��T�^Yw8����F���n�V�xJw�\�#ia�!��֪**y�����c��GG����P�����{����k����{8'�`�I\RXXh�VO��K
Y���ZzZZ99���~L\��S�� Uhiie��=:��?Cy�~�4�Ӣ"Y�m��a=W�w�˥D%�Õt���3k�T|����_Y���ϊ��|����N��0���N�Ź>y��#��6��@L�f�s$!f��ݵ���/��U�s6gk�*Xs��i6��HyN�/�V�*?���|��J���s$o^�:�)�&б��kE������:y�]{��~��'=���\�Q|=��P*=�(ET�h9��z��/_A-��k�(Ű���MU��� +��srϮH�'�+Ԓ�'�|��w�����"���B��,����]IM-n`pp��i��p:����;��uuĎ|�a0�w;�'�@����V��#Ot����N~�:�co1�T ��v�y��6o#	��2�����Yh�>�HƤڸ��g��~ k�߭8���օ�h�y=ޥd襃��8q��@���*���)�gDuM�gǵu++4�GZ�f;�hhM�B]TX+����;�d\
�dʹk�6���nojv�R�v�O�S�?�3��QT�����h0''�|�dUUU�|���$A���ԁ(VTV^�;tu�iG޻y���F]\<HK[{@��6���+��;i0Ln��}�߆.��uv*�����~�
}-;;�j~~>p�/{��f�ߺ����\�بkee养
�[.�<ј=q�m���������/G�w%⭹�P��M�5Q�/l�X��#�J/�v���,=9R��ib��!�ŏ0�0�U��JY"�ԯW1y�d�>��r���~�A�}}� KQ����Y�'�Qf�*� ��`�U�LN{�i,TN�IkUH�2�����vzb�	&�D�ț�$'k囿u���M*��P�$�@�a-o�曌ʯ�:�̣�W�^�� 5���t�ӌsxuU������`+�����������ϕi�����џ>-;�_�U��"�/=0�]��(��HK6N�d��o��;�)AK�<��C?$�����J?���x��7�Y�9���`�7�2���k��T��:!���p!Q	I�U�h����~r��=ǵp�GJ���%��C��%TE�5�/S�=�|Z��e�s;Ҧ�Hr��̇-=�#�; ��T�=St;�Z5�w6���M�}ֻb/	p�=��1���FryA�eGr�b%�57`�������mq�����^�����h���I#ř�e�Z��J��YT���h�ݛ7�P܏�n���͚y��B����z	c��=r�z��	���������<a��'�;��?os�-Ey	��K>�o�L�K���K����}j����s����}jR�#��ӕ������7{��0!�|Y�����:,��8���!��0���$�)��'�2+7�V^��O�n��%If��� 3���,0j0TtlBƅ�c:ӷ}��?J�$��%���je����Plll(� ��:��.����:��������kЦ�u�U�k���-��ۓ�����C
 �Z��"ľn�O�s�~�^�2�pӼ
�O�L�ی�Ì�"����F�1�m9��洳�j��&�)��o����[3���D�[�gՒ�i��9|+�k�%�@l�OcM�j^۔n;����3 L��k��F"?U� �ί�@w���Zyv�L�蝖x��2�g`p��:�~(q@M=ë�Ǆ]��*�܅ׄ$S޾B��yC��o�`�)���`��Kr�ժ'��_�U"�ȅ�J{��;�����@��/%� "��X����߅~���1���C�hħ�{Tz��9p�ӳ��ԫ��v�E2�����^����O�E�T�1�g:�8P	:QQ��՝$�����χ���ᆒ휮�#����M|��4;�P��ql��� Jߊ�1����ŴK���Z��W�0�5�Q�A��U�YS��H/�(�?p,��8��;�c�95�u���4���0t����W��E3��Vc�1�Vw$�k>��6%�m�u�t�*@�h;�I襖ʮ�v��XdC�Y�� YlQRV7�W�Cw5u;9-�'�@u������+]F���T�]���.�g�/�9`{�][^.E�C'�֟n�`���eJ(x�5��my�K=��4�T���	G�k��Fi�QtX���nLttօ�7�q���s��ɼ�f��G�D�ꂅ��"��6~u/�忲�u~�|��������� ��'�5���K�F
�����F��S��)��5Yf�0�P�ȦQ[K�<���h��a��3���~@7�)hI�
j�DMq�����	�K#�(���^֖���R��{���I�Y���}K V��+7\��:cMe-��(�����p�N��Y~׈�d���$�E�a�*z0��SnFT���@¯܍J2��K-�O� Y,E�k�x���x&aK0���׃4Z|, �F���x#/��y�_.cʣ�:yc���zT.Y�����ʧ��+W�{��g?�Y�6�p����޺�%�X<]A察��gT�Q9���3�.��W=�6lI�<o��`�[qc����:��f�K\P�����#�S���ėYl�gF ��	nR��M���ɷ�m5Z�r�o��r�Ef�@�6�ֽ���Z{m��2r{�WV����ڊ��| "��o��e�K4#���6�V�˝�c�r����B&ԃ���vP�����@)�h�#���n�r� �p/��9��w����O.���Ύ�M��#/��r�d#�-����ΡB�L�}���D4� ����R ds�އ>�7Rz��03B���Z��U����3Sl���1�$ŊD<zhp{p&���\2���[�v�G*]�uϔZO��*}�Y�8NJ9H���ў��y
ľ�����{GE��S��k�~eL�̈���0�L��i�(��.�V�I��0���h���6� 	�����.V�⵭YܼR��=^�8`f�z;���\��N[���,��p�Ü����B�]�����2D�S_�E�?�6P/<npM��6/��a���zU0D`b�'vͦ`�Ѭ�3|~��U��T�������KM��C0��b��ݟ Ȁ�iU�+=�,l(�%�w�����d�Ms�rtl�4�Ga;i���#�R'�4yǉ��j�����ju@M~���H�֬��`�U�z�h�P��W#V��Wr����}�~"|��yA�-EŮj��S��oj����9�����i��M6d~K�6�g+��>}X��Ț�J�o�zw[���p�ЦHBP���68M�:�������dc0�뉳���;�7�f
���y�_3�6Z���;�xA�$�?�"W9�HB��廇��Zk��"�� �r"߅����AAK�vjQ:����?���/v�IJ�Q�����j���R��辕Pb�J�?X	�J�&&���k��q�6�3s��l���/�i�+«�.�{�x��b:��=���y�)[�J��n�%�@���Z��R�w�Ǯ7�7L_��I�+�9m*f��7nh�+Ι���d�Q��l��G�Fg./pE�����l?^f��$���M2���F��Gb�rIS�T��Z���� @y�{��mݐg^�h6���M�=�`����yI�u�h��n�4�l9��h�����V��x��ba��Z��:�V�f_�����c��p{�y�Z>�Z/���Uj�>�Q+=v?[�V}r\�@���"
�Ҵs?տ[$�,�	c��~�+��ٱ�|y�WD	������`����<��:)��f����?Y�>3�����S��9asuƄ�!j�s����`��m[�>$���ю��u/JV n|��p6?���j��0Q�8f_ߞT���2l��.�7�@9d�V\�>��g	�9! �-x�eo�Ւ��P��v�Ϥ�L��cu�����hH��x��7��J�Z�/�_�/��v��Kth�{�%�f�<�H8�4�zgů�H���T�3�J����I/7+@ 5� �b�t���y��4�p���R�pU�#����10xAt�pI��Ҧ� iB���F�x�$�n����H����&4��������Dg����E�f�l
.�:}��\yۖ0�F�e�>2�J_*5/FQ�@i�&�QX�[�沩��'�}5��U�I���![Gu{��������&��l�������V!�qu]c��A�3�\����LM�s��|�~毚��;װJ��LtT�����^ UQ
��Kv-N�kX�\����f�� CC���U�ݧ��=���tQ'IMr�P�;$��oE��!7��#�h4�kP!]�R�/��� �b�k���D	i�6^����9	u�r�ʜq2DLpz?�~% k���,��j�]�����utc�	.�x�[g�v�4z��w�ˬQ�t���5�t�$(FAk�׼����8�7���t���̘b魎�� ��,Op���IdmDtoO�9�����O�FJ��[��<I�T蜗�.b����5�S�Z3�C�C�>Zj$���H �Ԣ9��E�����O�J�K���ԭ�b9��=,-Y!R�v�V�*��yb�3#m��Pr~���E$�������
�ʗ0,Px�` ��q�S4���W����T���;;w��4Ζ�6)�vt��U�]"�W�S�U}���S8��t�K���GK���>! �?w�9��k�����*��7�k?T����kIv�NH��x���*i4���2�J��I���|4R�����SJ��k���v��nt�U][�g�07e��Z�U��^�x�J*2�+#֯;A�)&g֕��{$�@0���ô�Ù����{%
�hg��)�J��$!ܸ�V�n���NחKͳ,;7��Re��?u\6: �3���j.,��
����A��X�7)��#��g ��;v�p�3_&3n�`s��1�,�nn�D�K��|,��8X ��|r�8FY��aj���Hq�)�$ĺWmڳ�B��6�*�=�	؀�>�������9$7�X`.`1�5�Ux�Ԕ��M���o�:�}�2� v�R/T�r����۸g��h H+���zV������	���uk��F�^(����Y� �N4�?���=@<��l*�ɧq���4z��F,lu�&�������i�]� ��C&�F�pT]���W4s�zZ��׸��q��N�v�lú���F���ʅ�W<���<D족f��[t�҈z��1��W�����%�7�S^�]���y=Y�և�ZsX��gl�K�7�-�{��Lt�gZ5�E 򳍍����h��Ϡ-��L�:f��s"��_�<����Ll�����8�ׅ>=0�5��"U�r�@�7^���aC��(t�K*y�Q�x��.��N �����E���j�@j�N��5�)�M&�@J�M����<3m���~������bbh�q��dQl��J��厡8���%�)�<�I<HՏ��������$Y8ϱg��r-�/�(&�
��~�L��gS�O
*$�+���eAd�����gc�zݺeP5�����)G$!���~��M.5��&G�I�5��{n���{>�\E�G!���U�U
�&�`�AR��-JOd�a�jh�$T����ב��厙f��"�+M�a��.����� ��WK�/�&�3�?�l˴�KQ@��]�tzMI� Cg kX���$�8.g�؜�R���-����D)=%��H*�QQQ��-� ���*YKO�[E�N\߹ůF6b�A�7��豹<���E\���t�(���y�Y�)U��j4,�)Ԯ�݂'ʰf��ĐVy��a������GO1�SC�!F��"P�������~��î�����'�k�5���_8���V"�/��:��9	���7T+5�a�.��5�W�z���e�� X���:�K%S*��$7���"aAab�����<�%+��"���s���*���m�G�iw"?�,<Pj��~�W#X��g+�Hym�"��;�&;jl��F�(�\�ҥVw���
�乻�z���8�������dҺ��TW�y��I������=�7��-pA�a�� y|���
'���=�<�=��Ap��$?���������e�!N▜ץG��wb�T�z��35���	��c.s��^>�@3��avG�(_�:�(�J����H�ǋ"��3t����S䃀�����K��} �
̠�}?ac7j��Pw��/�t��1�u�Z�x�&�8�0	ƗF�/%������M��J�U��jñ�Q`��M����l���黷�vԬ��'�>;~g�h�˛:~?me|�˴���̞�لN������&��{����K-�p������q��E`�Mє�ab/ ���0k&���.���s�	�9ТK�ȍ�� �N��v�nQ(ȞB����S1꿒�yAH�/���N�!�C�U��E˃�`�>�Ai`ńDx���<J�/�ږ�^1�f�<)i�l��`���J�o3�T��j*�0�S�z����hv��)G>U�/OK�C��$4�ǂT����9e;|G�sY�b�MY�N��"�G�eY��@�#?�����3�╲�鉍��p>@;�>�?e�y�A(� 6�hr����)9z܌�V����c9�����R;W����i���p�@C����I4�b-;cW��M>_�y@c�g�H�x�b�4oP��#ߎ�����{��Cf����Փ��?»`܎M"-G@���kT�ƌ�"��� 6���K"��ι�����lKQ�$M��������������L�Z�
g�c��1bC�Xڈ�ΘB�:S-��"�}���y� X@K����y$����SX��@�ēu�A�X�	Z�B��)�\���?��l��S�������3e_����Ú_mx����H)]d�T.s��D4B��ɗc9��< 6)��?�,]�ZP��l�
�y߸�m����A�� ̀��Gr0�a5���#[���4�?����qH��I��L�-#��Z%�a2�w\�%��*ۊ_{�~�TQ�h���pDa{ �H�U�R L� ������꿲�jS�uxq�:�ul�3n\ž����Ti�
^�d�4���&��밼'e?齸lK��2��CL�׭��dڦp� )IɁ��������Z3PK����D�5��Ŧ{ip��7��S|Vd�0 ���'EPa�<�e��b�����A�0�Q�Z�������҇�r�`���������N�vf�6U!2��7Y����DJ[?�ww�2� �{#��)K׼V�&�o�0�S��D�g�Z�nc֩4�b����~N���_�J�~����ߔ��V���dZ�g���x��Af�Ў�;Ku�j���"���ګ�2��̳6g�Y4���S�P��s�0��Ŕ������WLH�`Jnʁè����#棯�`C�W�6Z�Εgп
����1�sЗ�%��In�y[�^ǹU��O��P���FJO�R�[��O~�U���p�A���P����#F�:�`��+5O��f��g�᧑I�i��� �cIu��ۢ��W�/�ð�c�.[]6b����>، r���*�l�S	�]�
�4�;����]S]��G�{�b�ޗk�O�	��>'`��+�L�T�d�
,&�&����`�q%����I�`�eY��V�������Sq8��t�n��wu�J�B6���Ө|+	:+'�}��o9C/�{�U��cA �]2e�!���d�宝�_���lIU)��ܓn�4�>��/k%yr�,�I ԍ]U�J��.OJ��O����7�2;$�����,�R���\c���{Ū�~�MH �+y^)���h��8�6.}�'�ݼ�,�����f�i�����#��G����;�Hʦ�6����B��w�{8�q�Z+�(W�ڷ,�ð}Gas��t���(��
6D+o�㳢Ξ�-5p��o	�#� mܔX�.z�6Gh}Ʃ?���F�߽ٶ_�aن��O)�W���%�̈́���M�H�.I�'Oa��ɭ���߃)�q�֣�8�ttϧ_ ��R�3��C ���+b���zj���u/�A@���џ�y���ҡ�u��>�,!��X�b0��>j�q>�����';�q��{� �a�
L���W����D+ye��J�^�%�&dԲ����pE4R�#�l��L^�FE��	C��vg��O	����o�(���P������p������ �N�S���w�랇�)B����{�,����}[�4Ö>��y�]>��1�����=��K۟qd�Y2��R���i&㤅!���yǻj�ŏ5Mp͆�D��Ͽu�|���sL�Lβ*-����΃l����!)P?����<�O�kn���3>xL�)W�ɖy%-B�0�	��wF�H���2�3�.'�=���q@ގ�d��l���[${����h3G =Y�a����0�\�`�d��e����wMy[���(��k>�(r�|�J9&�����k%���S���/�]t/N�
�����ax$��X�[b/�E@x��q��y~�x���)k~l��K�H�j�IXϫ!k�Ay��_�b#R�B����嬡3'�`Δ$rO��� n	2�Սf��T7|Rp_�^�ț9�j����e	�)1�d�|���m� f�������7gI�K6��%��jC[&�|��[!/q�� �JC��+�M��mu����+��&���أG	��Yz����fɏQb����.|�M̬��}��6�R�͖�uڸ5��8�Xed��l�UKRҲ#�$�@� �<��h�fS;<�����	
^�j��L�Z.Br����#�U��;����5�XT�ޛP�)r�	��y�;qC0��e��̪6_G���[G�ǀ���Ӽ��VJv���U�s�j�^N�h~��u �V��{�>E�؞�{@]�g
�2�^���bN5��q)A��� �v(n�(�U���wO�I�sɸ',h�<_Yy9�e�^�`��h��r�.5k�g'!��i���#�xƈau����w���]#^�mI�9�Ȓ�}lZQ>�B�tu����H��H�_݇��ә�L��x����s��!$���X�|݆�Q��^�q�&��9QD���]0/��ff�<N��D�Y%� �'�W(2�#��^�b�>�����fh���ȗr�Z��ޓ�nu=k�߫����s����siP��|�/�˥��9���G�RȚ0���ѾL �s��=���eS����ۿ���>��|�D]�d+cy232�2�6�BV�^�Ql�[L���X�>N�C\*IV�<�@�_Gn�$�\�Ǥ������� �o�٧�����1������I�x�
�t�k��`ro�L[ʩR��C�)3��Su3zp6n�@G��$H)��U6x該Y:,gR���W���`�����@��G����).�����A$Qq1φ�J���B�A�keV��� �a��+���h4��Ie��9j��j��[r�}u����\+�D�x���>qFnO�J	@�s=�� ��x|[RNI-gu����wcw<~�iJ��Y4�?�4�`��dV<N���Ɗ�pw��&��Q-�y��i�x���q���������G%ݛd�fO��Z��zi9�z`�Wo���� �(�� �W�4�V��;���T���[D�����AAa��{��{���f�]K��g��~���w�K�L�5����k��g9* ..�Q-�즞'o ��2��>0�F5'��9��Y�.���������]��7_����?Xv�ށ��`hY�_��{�?�J�,���rL���y&t��s
�3��j��I�\iu��B�����2��Z9bBuk��G}3�L�a	=�Lـ���G�p���jo\��$|�>H�� o爩��� �����sH=T%��X��כ�w��z�01�>���{��<�j��!k�Lc?L1�.L�ʝ�J�)�<���zG�#�b��,{T �ssG���#�`^�sz��ҭ���{��-%�B���z�^3s��w/UzWpp�Ԇ����]�BpH���A�3q7���}S,E����q/zR���Qb�;Y����%oI���C����փǎI\"��j�{Tn�q�@	�ͳ��\K�m�T5�D'���Y���C�0���h��cU���^TF��i�[M��x&���a�����Ý�>�׬X�:nH�N�瞎����M��Q.����KV�{PdŃ/Ӹ	�5T��nߛ
��d#w�����������u�P�:@��b�6C^�-����;��?SJ9��_��M$�	1�5O«Ȝ!�I��ř�"w��6 �����6�>���*� X�,�hs%�� U�$��$���E] P:Ճ��T�FZ��+����4�,���>*�a�s���!4e�}'��ԿJ��Q`�A*�y>�6���%��7�"_@-�:�cJ
��f���1)�Y
#��������>��<�+3{y�o;�2>&����i���ս=
P`�-�3�qh�P� �i�R�V���Ǎ�:��wD��v�9��2���#wd���ڒ=���h&�b��Ёg�=�L�k'O��Z�)�� K�Y�dWxI�M!$_��x���c̔��_��Kc2�a���lˡ�?�ڒbԂ�u3\�X�M�j&[����+��S��ގl{�����u��骧��!N�-㷙���sN�{e��� �ڢ��7�dV��/Y����!'G �=��m?��V�<�J��Ӵ
<m���ω=�������!Eg�:v->}O�u��	2`�����ďI�5��u\�U���"���H��2�7[�A9�:�U���+�|�u�6�cVmb��o'j؞;�K��5����:S��ȃ�/�����^լ-�~z[Y�k�I��gV��} �{��8O� ��`?;�cI�9G1�����/&?�`�l4���W��f�-)��ZMf��^e�!�y�58DC�'q^S'��T\v3�0���B�Z�k;���x�y5�韼�DY}�V��2�j|�+�?�Z�:փ�?& �	@s��s����Ȍ Ypg ���,�f-$1aXaWs��1>�݄�$�-�����Lk9��r] |�#�f��sM�:gUo;\�
��3�0��������5�kҿœ8�� ��A���Mc��e'KdOFB�/���s�U��Ђ�v��j�	��ǾS;��?&��xཀྵ���#�x��[W���\�r��#���~a����贑gl�
��~#���
���r]�[Pt2b��57�F�W�fs��t��X������FR=~�n9rc��N�0��Z��]]/��S믤�u���㷭�jmltl{$��śH�m�����8�9g̃.P�N��>�ܓ3O� P��F��x� Ӣ뛐\Zrq�K����]^�lDP�ڹܨ���Y�Q��I��3lh6/��׼��	*��SV�%���S���t��1ۥoa����Izp#��^���M�RHV�l§S��hHxc�ໟW^v;�0��D?y�Q��m6�2�kf�Q��{$�/�!��0��(��Z�k?�m��;�p�V�=�x����% E�g�DP�S�fo$�)���b�}܀�ۨ��u����Y���x�Zj�4uAj�������d���Y��#'�6h�,�cݜ���$DU�/݁�>F�����R�q�����][��KW��s�5����$�VI���Уm[i���
XCa�/��U�mRL�&%�^�N��'�(;��>߅�#�d���j��v��_랻ל��P\zBjx%��=��a̹�;n
2�x��/t�A�Ң��z��̿}� �� �'r[ȸ"-��j��%+�TW�6B�׌�an�W�ٗ���'�x����e��M�/�p�N2u�&���) �3q�Z�!-/v��b9q)nxXW���Վ�s��X� ���������dT�Y��?��� ��¢��5�!�R����M�J�X>�
 �x=�Z;c�f�䍙�j��-��
�E3��Bm����S�!����ͧj��߰��.�zj�'�V���z{�#^&�b��d�>qȋ��㊩��L�ΛS>]�}�F�	� X�u��i�x*���VL��������-�`���4Ot�*.S�޹�,�@�eL���V��Q���v`����E���o��7)���!.�n`�� �5�Vw/Tb��m%�����S��u6{�
��k��2�~_鄏U�x�C��=��C������D3.Y����|q�p����E$y7?�C�d�F��W�����b�?��E9�BG�l�wJ|:M�����yT��[6̫C=�o޶,�����D��s���w.L��l Owٓ�Q�`��V�7E�}��_�DO�|��j��$JJ�Bh"��_?B�����؍��[+)���KR�60e�ڙ1r��)a������⧳���R�b�˸r�3�������Qm��CO
 �rk���F{�1�V�M]_go:����������������� 2l��Hy�e�\�9���|��H�X|!c�<kV��VN<��B�p�5��MpQC�e-ҽI]� C��.70 ���_���i?+6�����-���<��j�־�\G�;���Z'xgF�Ԣ��IK�����[}���F��ڐ".����r�A졉���h�}bYX�w���p�p]f��w$[}����1	��vWߣ��;ր*��k��+�����d(�w���V��ئ�X��Uq��i��8)b�}k�BY�L"��@38��0�3t(9��1<.e�u��ʛ�0��T^V�J��,I���v�����S��H����H
k��޵D�k�#Eǐ�Do8!<p�ũ���ٵT��/I,s#_&s���<����I�.l1��� �j/Cq�ֈ���-�/t�I��?�Xm/-^릭r�Koٮ���-C��W)�)�6�H�_l���hnq�=||���Ǘ�2S����,�e�J��-p���O����\��8US��Sv�_;���O,(^Z=i�=�}��b�����".d�jt�٪�[� ��	���������y����z�J��\���'Sa������;��\7��Ȱ_%!�t�w�B���O4SM�N�� �\��9��W�HV���OM���K�\��a��ė���x��pʆ![�%�:����?d����1< T��T4��3�)ۡn�P���>5�|^�p��@⬨�4������4�3�2�~��_�˯ztn��b�n�X�F��g�����K�<�8e�F򵓚<��b��鸿��*��9��5���+���M�L���l���ݖG��G,�h�������7��#��Pw;Q9��
:Z(k��ͻ()z��c�y���䝩�T� 7y,�_x�|J��קѺ�H�ݸ����6)	����hi�2b	�,,��Fԭ�NWx�^IwV�&����*��I�֐��V��DE�����ǒ�O�^�ޭ��i���Vɗ���L_��j��oy��׌�8�����k�K���JJЙuc�j� 9Q�O�V��0B��x,����lt(��j4�$���B@]�JԞ�v���y^�EW#S[�.uW�j�%\����p��\l՚/2.|��V�wf=֚� �eG��Aǖ����6�1x��ML��u%*Ѷ�)geVe�eQ�XF�%r0��K���zi��a7~��Ϫ����6̞���w� i�Frw�L~���(e�q�7|n_��[���ɡ���e���a�Hš��,]�Æpe��kjVT ��ӈ�Ǵ�Jd���x��|֊��uUuF�v�3���c���^N�Io��S3����=�G�����C� �����t������-�X�a�"�����B�������[<g˔F�Z�%�"��/	W�e��<�g=���O���)�˗bG��DL7V�i���G8���3�h&�����}*ɞӧs�]�ItA���,�����he�3~�r�>7����Z7��.o��Pm��j��UҪ�*Zp����O�Ӿ���y�v��cI64H�g�e`����F�LC�Փ
Êн"_]�W���I�j��4��j5(���}��S{��̙Tsl�����r�$�C=���+4�,RF%~�g����:,�uR�MHjҖL$�ڐOV��G�Z�76J���-�l�[e�c�l��f�j�����5ˉ\�[4<���y�t]��Ë5!�$r��ߥqw�
$��щ��]� �!y&�����Xl����V�B�ن�����;�B��\����yA����i��v�T��xGz�:�$@�(3�,���GV>w�FXk��� �瑮Y�-ѻ�B����ڶ�J���]F��k[��K��a%�t܍�B��D��,4"�r5��K�G�:k�P�cU������X:.�;O�ט
ڒ���a�����~<fbA��X[�w4��`���&Q�O���l����H.g��^5��?p�w=)��vU������}��*]t���_O�I����d7���VK�q��	G&�}�����eJ�3N�x[�Ζ�A�<fe��R�2���r�5�s�����d�-��DI�T6P袣JYբ��fIz�����r�rz(?�wE�������C�W v����l�W� �n��M&
����҅���Y%��>9�)��㮪�wx;g����ȷ��}�����a��M���ಊq/�����8���o�ļ�g��q5������^W�i�T�̆ њ*Y�Mp�?�x�aXb�3�ho:ju�=�C�ʲ}߬k�e�"7g��t�C�3�4��'Μ�)���Mo�鴡��7�@٭��u������l�f�C���mr��ӥeÚ���w&+��k;�7�yM6fn�O�_�4�i�/��_�1G����/�@w�xa�7���)�u��f��|G��y�%U�np�L�k+���~/ؿ���=3�8.;����+qI��a	ʻ��KQ��$��Z�1YM��}��×N2�u5O�L�_�ļ�J�w����-_�ua��$�\l(+�LT������+�cmQ�"�M0��ђ�1)��h;7�o���$�?�@�E@�4)����?	Ku�ϖ��Q��;�Z\ibW���sV{�)�C��`�X��M\	���zM���r^`��;Pkȴ'�r#W���).������5�'�T��\�7_��Wh�J7OGdK�Y�ȮᕨY��X9����	I�Z�aiSF�Rړ���]��s�F�&��B#t������k+xj�A\(l��>�JEe>K�w�DQ�����M�yo�������/Lk�֌���?����ؑM�Ԙ:]sӏۖ��Y�ܽN�E�����C���]�����G����\�
7�MǇ��,�8�ȟa���a�ݬrt�j�rJ�/�8)M5����C�=V�0�(��X���ߞ�.U"/V��tV�C��=��H׊�0�N"Bdsja0�+ETX���.�Q5i��°�v�ˋ��ߒSe_�\�g]Y妛M93��9��់`�B1Ӎ/])��|�+LT)�m����E(F�X�<f�B�c��KB����(���n>,!Ry��P�
�
dH���f�i�~R����d9X��A!'��*vR&д(&�Q��U�to*D�<+�<�W���)%�h%,����ܻ��}F#;���Ĥ� 	Uc���Y��Q�����@��Zv����usb���cw�b5�PW�Tz]X@#� ���r����T=��Z�,��j�9MF�}�+�xe��ӵc��/J��\�QW/�2_�l�c����U�+jXh �i�ݵ�����%l�vW5VN�zg��	���1��N6�? �
����P��dǲ���c�62���Q�F�X]B�|�F�G\-W�5�`�V��a5X�p�p'J�~�*�bإX�֔M	���{*D�-�Lߗ���5���i6��e������g��q��0%ɡ#\�����ٓj���F�Zl���U��f (y3�2'��Պ����_6\}�#�Nѡ�ϙy�F	Q4.t�Ӧ��Fp����c_bɗ��3K��k�ZЂ��o@�
s��^ۖb����e�K��H�0(��;�8������T�u�#/��޾HS��[�f���0��'բ\̓Sǿ:��ػ�M[��X/�O�Y}d�ٓ~��̕y?���C�bV�@>x�ι ���%��c�z�~A�>>O���Қ1�.忒�o����P}��Jl�{}ե�jp-����D Sx�C����>�t�U��`���z�Z�_�+��� �󪳩Be4��\��ol�|Oʞ�ܧz���/#f����K58��!Z��^ᤑ������~��h���K�@��υ���!�������˧��E$&}��FM��y�\�x3jnݲf~ej�V汀t-��>�}����P��M�77�S_7}�3* �ؕ�����7�q���v�/��H��%~7���ԅ�90�.n�:c�ds	VAM�L>Ɓ��Ŵ3����sunof}x=��J���1I)����+l0���"�O�P��/.�$�^5����<� ��ȳ���`��Ԧ./6��eL���i����ơ��.͔8�f!���x�Y�a�n�>�SFy�����N�������L�|��&��'���c_�6 �&�k1�pև���a�KⒶ��+�kr 8�*9t$�BP��^"@�)<�{>�������Q@Gɗ/�D����a�$ �y�Bs�A����ᯟ�-K�}&_E���������Hχ	_�n�q�'�B���B������濾]�\S���7v��(6,o�H-X�{�	t���͵�ؔ�t���d&���c�A� Jiͨ�ɗ*^�>��[yI1���4�D E'�����ڔ2Ta+�R�L���Kf����̣�4�1����nh?���a	\wF,v���8Bd�ˁq�y~׋�/ {�7�M!M�	,lJ�Ǽq����s��H�g����C�yx}1tMS@�.��!U��/W�ڃ"SR+hqh^;���/����ӕP�5GgE=���Ի`ݒ��v��t��"�c"�51OB�&`��/������йu����L�rxWΑ��/CgӄC����MX��i�%�?Xw��xj�w�j�t�-n��.	̒+/�Q.�'瑌E����o�
�Yq#�B��xy~�0�� yn�g΀�PQ���X�{��L7XT]R�e� ]:�E� ���ڞ�&�+���H3kVX����/�
��iBO �oS>&��><�rL%g�-�{�݄m
�n�7ۼ�4VK|&v�W������3��;0}����V�F��^����ӛ��i���7}0F0d�=_E&@��7ł�,]�]��lH��\Ј��(b��b��f�+��;w�Z��J�D��i�m$=��s̑Q�C���yh�}N��'�����c���C� | �	eA�����ε���tǖ���"�ڴ{]��V}��O#>Ȉ A*��x�U\Q�q���+������J�a�-����nғXuZf���스1Cmxh9�����jL@*�)�����&�(o^���5��4�U�:��DKu�g��`3{�Hf���q ~��B����|��P��*�rW��R�S>��O�k?���D�1~�v�������<!;�f�9x�^�nG��c��)�C�Q��e�P���|����T ?��m�h��$�|��s�ϒVkމ4�,�]�Eс_2=߷B�~뫄N熫~�c��*Jv;6E�;�Q��9ru�c�.i��DG�>�oJ�_	V�FҚ�3y �:�p�>�-��G�80X��)�>�\}}��r����jw�|����K ��7:'B�4�N��0��b���C��2�Es_$��Ze�
cO�f�:�;���Nl;9?K�1���Fs�l��>V-�!����L�a��,@,�vN���ɝ-�N���mcGF�\��r*X���n�[�<F�'�%-P�9��[[��[�@5Y��d�Ł]f���>ǵ���оB�����؇�%F^�t�&�)1]ܐM�*4Rw���X��t���S���S�#����?�o
����{����^��k���`�m-'�d��_
md�`RJ1�.<�<^���R@�Vm�vБ�1�!�F�#���M���uYN �E�����	����tj_1�:f�KS��iW�Α����_�BXN���A^1)+�ޅ-�?d��<����i�2T���)اί�����6��yR��7��3Z
�9�	�5x9i�J�8.@�d�L���|rʐ%�G����O��iZ���^a�0i�:|ްt��/*�;c��[�"tT ���/J�����Y�@H���+=�<ŨMm�@75aͅ��
�i
��M.`�SjSٚ�q��8�n����Zz����y�Ou�t�H��'�&�B��a���d%��A�5 E򿩿	1�N�Q]��ҕ�dͲ��<���{FV����22<("�\�hH��_�ȋ�L���.���,撿=d;�.U�&N�I�	��R���eTw������D��M�,���w��ĵp��[���/� ��-@Ҝ,���(d�r��>���mc;Kv�Q��3=�J�)@B�h6>��C�/l�a�OC�jpv_�J�A���?S��C�YC�:JP@���T;���2�~����s�0�S�+J�����֥�.wVU)�q�=���7w�1�Ώ7[��1a�Γ׎=a�<���g��!�V3k�c[��c�7�Y�;Ĩʦ�偩%̏�,����$���ԇ^FQ�$)yV���e�����g.��\h�V�߾���d�KS�.�i��w �X�lb!U�R�1l#��ݺQ�ݬ���=%����s�F��ܣ����s�F�P˔�k��=֬��ϭ6�G��4
�h��5��B���� ߔ.w�!�[X���MN�S���iG:�I�p��`�cn�݂$g0
���������5�$���E�$�&���D%��К拿s�& w���5*��j�-�K��J����G�RҒx���O���H�!$X�I��t��h/����}���k�fژ����)����Cc�i²���� �߯f�!ȵ���ݱ����]����Gj%�5:�ix�������gC����6.�dZ��~�x�2E.�T,��Uep���/7oH�!�tf��T9z�N�=/.L-���F��|x�he�i�ӎ�T��\rK��L�狳�5�M_ą�^$ؓ�.Gy���=/�W.,������w�������b�K�:�Ug&k�ok�Xfn�Y(��Ӳa����
��+c�X��:�6:w���p�E�b̢��w��Lŷq-fZ�vn�>J@��2@}�	�4m�Η�@�����;oD)�1Ԏ�O�P��?�ک�5Zd`�Y�-�K��������*a)RA١������:�o��=�O�3n��5�&�vh�ٕ<��-o��G#L��8 %sљT�Ցu*���z��O��+��(�r��Vq%�i��#p��f�_4�wn��� ��p�c�c&��:� AP( K9p�����a]�	�1a9#�ze&s�
!S��}��eP�����4T\\�jťƤ�>�Ǳ�b�,/-Hp@Z*�$�;�m$�����՗����j5�};�������u�F���[��4�lz�O��e�c����	�D � �^�l���jG?���!��+ݼ�z�R4���|$E*��@��W$U5*|󿭺�Ӣ�V��;/�NN��y")P�����dCԄ�*bF�����j��,-���8_�������^Yf�O����!��1�rX.�xo��'(Z��Bi��Z;�G"'޵R㺋&|��m,�I|QO�f2i(}쏕b<�oy_� ��@���i/��IPL�̥r��x%�)��k��U��R�]Ԝ��i4���b�e�@�ha(�}P%���CH,�\����J*v�.�
����4�j��Ƽ���4۳ϳWͨ�UĨ)Y��r�[W����0p�*���*��6be���@k��Ƌ��G��t��(8s�kզN6ן	��rW���jX�j������@�r+�^�qu��$y�����������i�UNm�GN�ú�E����F�ԕ�ǦC�T�v	Y�	�}�ݢ�і=�7F��?t���l�pk�g��<F��]O���v��> �N���@�-��|,T���:Ƀ-�4��w��a���/�v���J5����y�Lg���_?�,_d�d�VP�ü����ĮM-��LW!E����)B��#�Up�M�i9t����lI,-��k��T��t\92�g	0�i��*�dÃ�-ZU������FW{�;�%sX9j�腺����YR�>	o��m�9ɬ���E`�4e���(�x��%地`���G�!	\T9yv����!?�M]�������\{f�*Yj1�Ez���r���h[��&�$^��fG۱�y�Q���ǫ���xh��U1����X�Α�wm���7	�w,���ܧN�|E��Gy�s�2j�V6���/��kk��t�;C�6S�]���3G뺼i՝�T�j�.)����0�5�|B����Q)��y��V۫��H��ȾUZh+{]Z�Hǣ�T�R�\F<��t�I��M�흥��Y�;��XY�5��ۮ������yq��c���ZkX�K��<�5�]�n��� �$�`�G���Q	'�ms�=���H�S��*��p�!���c �Q��h��j���f���y�U�ֱ�;C��ڍm���V��jW�+����'ᵛL9�ڧQ���ŀpY?��[��
�o>>��un��7�c��>�]2/���LǗ��re��R�iRD��uk&���%��qY�s�&Y�����������%�<�����$�T��XM���l ��ګ	vړ⺸o���{T5�\.�6g�-�A�_��|��B� ش�h�'�Y��O�� SZƨ�@�M��f-.��[W����O���a�����2_F)�~}�����ܹĺ�b Yv������k�0���r��c;�vm�$��)������hn:E���xT�y� e,��?�[W�H��:M'����a�B������SH�{�.s�fEީ�IA�<�`z����ax��d\��%m[�KA_��m �pQ�>ƺ䓈H�D�:���R�|k�j)���YKk�ݨ�Z�Z F�+QpfGX��7�X�6v�9o�hP汍W�Vx&^�%}�f��-�<��>p���B.��?}pQ (B��kP��m^����B��x��!0�ѫ6�x��_�h�w��L��f����a<Jfl�~���w��ٲ@�1��z�!A��A��O�y��!��v(�"<�� �����c�̗�b�(��	:�c����}4��:u�Vĭ{O�%.PW�o����Xb
$:8t9,r5�;�L���P?��H��c��Ee��{c���T����"ڜq�,����敐���s�0�Bn����)��'����2�gk��>oV����B6��"?K�8�7�AY���Cא���S�nG�඘���V���^ѷXϴ��\Oq��RSb6��X���������)\�
}�Έ��r�����X1��/�����G��4w5�v8���k̜�`婛�Ƥ�����2��⼹$t1;�B8)T᪷�]��6gE|F�� ͂���G�k �$D�TE���X�N���#�ׅ������F�C���_��,_��2zi�#�Sh�?)����a�&b���Z��sU�ێ�a�d6G��0�|��J8	hG��Pu.<Џ~Q���"�u��TpW�L�x��Ȃ
�i�`�-8/�}s>_�^��U�i	��6*uNYi�-����\����w+�Yw PT\�������|���]��l�߅�hi�&�Ŧ;�ݟ3�\\�3�{W��C���m�ѩ�wD���"_P�)l��T?/uT	�"Bvj��"V��pv���ts�vk�#��C�����b��ܹ��z�����܄m��яg1�?#Lrd����Q>�Ypw�r6'�5D��w��Җ����
�,�;i���O�3qԤZ�ᓦZ#�C�q������:����/�n������Ғ-��7"��� ��t�D�q3�o���	���[uoP�]��E~�����z5ռ٭g嶓(��k�^&%��VG;i��p�8�ؿ�k#M���N%���㦲�'� J2�Xa��Hn��[V���J��搣*�����!�\��`\���:Y����5�
�����t#�%��J@e��r��d��}���]7���YiU�	d+��0i1V���\����s*��5�O�?��p�B�\۴q�jWV�����j��3���?�սC�o�_����'�[��؉$�ܖb!#�����顰^�<-L�s�Nʎm��m��ݵ�T��ǲ�''�;g�4x�ۡ�L�l�"�:@�J����6�N��@��P�������<O�Bk��gm�tm�a�Kn�f�m���r���>}GVC�}�JD�f�d�P��$g��\����+o#��<x\?0���|6�vј���ުަmb�$�)Γ���Z�vJ����]�Y� ^v�,�2R����q�"k�E���I��P���>����0����9[�lH|z-�
̬��@^�	��r=���K�Ŝ%3��\���*����@���+6=br�3�W�k��%�������L��`ak2ׄ��!�	�-���lHQ<?�Ɋ�o6��� p@Gu���_��B������#�W�U�:�YG�خ}���|2km6u~ۛ��ܟrR6�N6��SL�!�r��t�8�AN�����=�g�8��h� �ɾc����9
)�C��§��l���'��ە����PÃqV�o�E����ݧ}	$�&�>���o�<��]�dP�V�!Q�!`���*�Y�l�uɀ�I�uq�nn����5���w�K��I˨C�]?��`�%�G�6����!D�E��t^�z_�=Vɘ�m�3��g&�3�f���������������C��Sg���t���0��1}QG��0c��XX���d��� ��Ѣm_��ˑ����'�u�i���&`~��=D�?���涋�� y��ohgQ,ԡ��g��������}
m<~��.R�n�Ԓܒ�n�2�6�_��6�m�����h��X���QG��}&v{�^7���浓�T�L��K.�VL�ݹ����
E�!��k}�s��o�b�Xb��	~�ɨqk�b1ц��7�ɓ"^e��H��ƶ1�-�Ҥ�SE�a����< �%�LW�Qk1�D±XRP�{Y2�����~E����D(I`oi�����)]"���Z^c����_nF�����r������/������T��v�#�aʁ��ҷ��UwsG'��eT���<g�at�.��5���HxN���,L�d�
*�� �.v5�>����K֛I����m�R��
 �72��l�D��	6vSGe�f9����W�*S1�X��Z���q�oV.V˖�?�&�q��b��+:^��Q9�(D�[���Ϳ�r�;,e��%vh����RM�^�i����l�:��*�0"q�RX�	�zp�N?d0�e&mxG�a�۬��>�o�#�F��a�q�CZ6��t�h�m<�︋�d%_���&P���}���k�.�s�_A��?���ݱI�"N���'�?�	�tx1)+;)k33='�UG=�܆�c	����pnx !4�F���bg�Y�/�V�6�U��u�?7��lcG�*O(!k.5&�q�����9�\ZLI��N&�.�	�89�L6V>�˖���䨩(X�H�C���O���rɣkWd�X��i+M�K��N�f����ʩ�hw~Vo�kh<�(�����'s�GMea�nP�.^[[�$i�o�Ts�������.��m���_�Q�&��z|h@�%�c�v����0�5>��s=�!�⹡X*�$Ӡ���Q���e�v:������۱���BO��|>�~/���1�������(5{��g�l�_l���?�WB�n���9�5Pe�C�ǒ�}%���=��"C�(UzU[!�C��g\�t���f�d>oж+��Œ��&sl��:
{�]�,�W��f{�V=I`��3�` �l���-���j���h�2l�n76�ߧ��:p���d�υ�s6�q�Y��p��<�g䚕鵼7{|���MX@f��6��qr�����`�|?���>����Ә�?�O���)�E�"[��Dɧ�<�$�\��>� ��"�J9���.�o��)oZ���;PyЄ�F�7Zn~s���>��;��8Yf���;��uO��}o� 
&�q�ޑi�kO"�� |�SR�M��i;k/u9�.Z�
�+S���� ����r���~}��2Ci0���
����e��f��Nq$�pf�$�J�!ҳ\N�6���Ra�5���|S�U$�~�� 1�C)�����2|��]�%���R9SU���?ơ����lxr\�7�d��]/��_�����38�6*?6��P���8�xE�f�8w	��Rt_��\O�o�`H��x%D�b�p��7H�}V���R�p�C�r?-��[��.p�M?�)�Kr���d.[#5RnLԃ-v��8l��?\v�}Ab��B��k�כF����wG�"���4�TU(d�]&÷Q��WV> �,AT�;?{����\#3T������*nGa�4�L��UĚ8��E��bu��dՕ�4q}��*�W����[��
w�3$9I Pw*l3&$Db�д��YQ������PUM'M�	>�d�T��N������ڍ家�m�vZU|��h��k��������s6�@�0�v�k�(�� y�c����/X��mS�T`��O����~�כX�K��H<��H��i�*��i�(�i����M��'UnJv���#w e�{�Y�5�|j�����n�2��efL��ܟ_�]��o��N�q��H��u��IuH�_��|�݁�*�1n��iI��q!hu��ct��W�l[�s`��������[�гJ�=\�4�T�-AA�G�I`�[�����~�2`�"��N	�F5+b#`]>`�+��(^4;�Y�d���b��ee�v/'�3n�gms5���B����l����qN��lﯲ\��wUsu��@�K���	}9�Q���(�X���1�s�3�޾:����,㟿}Q�XE�w�^i�������6[���<�6�|sl��UCn�+t�����y�(w͙ctP����������?�F�Fw�"��Ϩ�?� %�
FWs���z��Y��[��:��/ʵf<8�ϱaկ!C�h>�4��T����*��N�1�U�J�c%�8T*w&b?~�����?�@݂O|�r�V��h�qNO�x���v�����朰}\�J)��Pܥ�e��Y�I��|�����B�i�x"d�z�w�gb�QN���q�5�4D����	�M�um>��~gTQ$ӆ�L�K }�,�=�5̏�UM�~�;�7ͳH�[2���U�S�3�}gݒre?�O+����aH2��-E���@¿y?_e!����~$,��5);�7w'�4X�\��:�t�S��(}���"e;I�,�t����咵�/��XzU.y�n:8�V�6�۳��V)0�6���K\�μ�H<��P��#A�PT��v�0�����s��c�^�@����_j��{��{��P��}�<���x�ap�>�ff�ӏA��4��Eë9=��;��Z�@��a�@���U����/xBy�T�f�������	? ���H.�_�u�[Z�ǜ�'\�V��:o)�WEW��uD�wi����΍&͂�v�ro�bP�G�)`�Ԯj|kc��svDu�u�<E��K5'lE�OՓ�T�����F�g��@�(�p��/�C����ԏ���]�Ӳ�	e����g�i�2p�|�"Vᓂ^��t���b�]��D�)1w�h�U?;�?�Y��VJ$`�v��}�U�����7WUe�dm�R�%�秂T��w�ԙ!�z�1or�����-��0�lC� 9�UW�|6��ǚ��@��DF��Y4��6���WQ����>0k^�5hK.J�>jw�]B�Nю�>�f?���z����<zG�5�F��M���4�߈}�_���ztz5~���+��CF��� e\z0�}�\�m\��e,��$9̏�s��_ۍ�h���=y-7�h߶��9w.��d�f��v,g�����;>����;��w~@�|���eo��+�sgq�9���*��&K${���e�4��C��������[�~�s�l�h�1����i6�#�o�:����.�{!�����`�[�!��xc�	�>��׳�	T+2}�1i<j>[z>�(I,������<
����Z�����79˟-��pw���/�p5_���ӆ�-���P�}�_k��Q��j5xЍ_"��T�1�T�b����*ϑhX�"����W-��{�ݿ�%Z� �41��;A�� �Pa[1Mw�DN��Ơ��i:�ru�%�}��<�a��<홇	���.̔���s%���������P� �My�����3�0�,��&s>��s�D�y�[��o V�����0���]����O��H��
��~gwf���4�dB�7�zq���@6�CY��]�#	{J���Yު��gO�k���;��O��{P�_	yj�E�ݩ8iT����{4���y����whg�XAR�s��s�@�˧�ssC��:���k��āF|�������
�(CT��HC_J����缇�^��k� ��;�7�o[,n�詘�ǈt?�aq�n"V�74C��*m`���a�������̰���0�m��9�q��?��;��r��'��y8j�X$^��@��b�9*��k.�f�3,��۵+>>SH���_l Rt�9w\�%rl�p�ju���Q�Y����g��j×�i����Y����p�ƴ[�Y1w����v1um.�pI���Eԫ�2�o��q�E3ī��D   5>���rl ��brY����Kt����ϥ���(U_R�rc��w�;<	e`�#�����3�E>����5�*�M6i�n���t�d����O�Nq�غ�@��3�&.��U�6��3�����x�.���� 9�E�^|Y�9^�>׺:�_�#��&b:˥����S�QByu�C�R�*B�����ziۄt.)� ���K���  ��t��tI# 
,JI)!�" ]"ݱ4�����y���qTv������ra
R���z}�/Tӑe��N�#�[o�ֿ||����١���?��z�zWd1b�Ջ�@�wK�t=�Ë���%ڃ�i�f	d����UN;���׼���.¬.V|>
v�;���~�>~�6-^��۪�0�,��޷���T��E4��}־<���6l�,��M�d�\�����W΂��29ml�[�g7fO�v��
*�N麭e2O}���_\��:��Ѻ�a��
=��7 ����`�|i�Q̶�+��`����ۻbf����{�~����"�{� ���K�$�.B����jXw4�:YY��)�tͲ��z3�Uj,��m��qz�%"�֗��x�V9&��"�To2� ;���d�YB"��PV���ɠU�h�=�F�lim���0])\�u�� �gZz�J�X����������n��^
���g�?kZץvͬ������
՛��<~F��^_�g�͟��[~�n��lQ�%u�������,��N��VE����w��˽������??�5�z�X�BK���w`�ef�g[���G���S�O�T��n]�F��h���ZMa����8���b�*=���r )��Qs��ec}ƾ�O�0���J�����2��)�`7�obg�W�Λܞ�~�I�O ����gn��r�x�ԡgg��CZ��*�o1˸|�+�V�XN8s�歘��7�S�E7H>Ov8Ϡ8�qHJ���5���Cv�8J=.��b˔1�fE�H��v�k/w��>,���Ŧ�8Q���0�F��Z�:��t=n�^7^��o.,F1�g ��y~�m���Bj.'g�|��>�+wR%8R��Ij0I�1�_np ��2��{4@����+
�	ؿ5�F�����[?�Ia�"��{TS4��fi���ٌ�ź@�j�ﲖ�݃󲻔t�U��NuIW�����C��$�/6F=c<��H0L��9+�1Ҫ�M��e�*��Z��.�d��O�RV�|�'|~�)�S����X�+���	�A�@�7t�h�g�G�團�����d� �t��^�nx3_�׽ay���е6����̴�����n�@���������,܅��,�r��%��� �a�6e7������s�#����Q�������=��7�hhU-�/z0���1����t*�y��7"�?rdU�
6%lʰ�I��㺎���]�e<p�¬T塾�����<ݮ
l�3?����yt��B���{�zoͮ�s��b�HDW�A�t��"�G˼���^^�hZR���5���/!����R���&��tF�v� ��d�%��?��u�T��R�s�g���WA#����~1P� K�h�����SB�xt���s)p#��"\���[�ܺ_u8F+ȁ����W���������vy����Xp4���lQR�����g�}/2�^9k�b�7�5���y� ��TR���~�oט���E�V��%���О���S߯�����o��o(.��P�:��L~�ӣ}���{Ճ`~v�_�S�O��\׮��Y�屼�qxa�q!���Q��ηッ�S�'�����ϐ7����{��)ݼ����)��*/��}A 5�###yi"���O�444�w�il10�K�J�G�G.�tl�I޿%$iH�A��$a�w�I�gB�M�e�9Z+T�X�ⅱ
Sf�x���~�=j��.s�U�����t�������㷪㈴��{�t�!��R�t�So/�O�Tp$w']N�|�G�1����W#���$C����ŀ����ME�WS����G�|�Y�[�<��}������FG�vww[��+���:G�z�A�°�T���=�����,��`�q)�u���U�t&����ۇ�(ޒ? ����&����4��#2*Wm��j
�WW�pt���)ьx�w^��W�&��o>��*��W��7�1�#�AlY��_0����&'��+J�[[O;:X�M���e�,֘[��n��se�Q	b(�
G����Ì�V��U��ߊk�g�A=�[Ε�1���ѺS4���p�0���K<N�������;��ۿ�ONm���\�jE���O�X2޸�B��@y�hz[|������f-G�^\\�����>���䖐��*Mnmi�655�'"�9��)����h��U���$$"�����{�X���M܄��N�J���l6�}	������y㱆�m��7^޵�M.z=W�^���^]�ϋ�[�%F�B��&��ţ���YG�2Ҋ�R>���;���J/��e�~\6���.�?'�-ύ��8��f��~b*��)vt��9�+Y��6�@��B�9��c���KH0455���I3G�LK�LJ�00�j��R���aT44�-�0M�����\�������Jh+*_��_�3V� ��e�S޺X{ځ��] �[#ܜ
��� ��q��*d!$(<��{v����G����v>4$&�㠎�݈�ř6b�K��y�R�e��Ku"G�'�4/[�m�e[���x7+�)���������?⇇݉5*RD"O��B
�	��d��o<��CYW�?�������F�Y�BfV�tth���g77�H�^�����o��E�B
;�m�����ĞO4�4�n�گ��nѧs���X��>VbR~Zy�'�w�A��%�46]1��W��JKgk��i�XX����|��qyz�:��Bj;���{��b��&��R�#-�aq���w}�=K۫?�W���-��q�C�-C8cdFG���(�^��������Y����*VNN���öJ������Ӏ����tq{�fw�;a\b�`���1#Af��8K�����ȯwX�[���8I��c*XM���R�g�1��ѝ�P�c��
fI#Vm����Y��-�F>B�k/E��ju`�c2�7���7�Kte������Ӈ��6�8�ﱮ3I5��H=�&���@tgq�3J	�������F}V��h|^�")ɨk���z���g�acoo�g�ںI���g�d�$Ȩ��Y��VV�)��k�C�&�AR�6�������:Z�->��SG/&�dD'�
�������X}�`e$A5"�oh�y�~�|�Bi��e�K��9+��uLp�e^��ܗ�/�H&�xܵy1��MS�Kn5������/Ok:Q�2�Cvv~�]
*��|(t�����H�_�k̎e����C."m�0Jw�33@M"v'��X�s�#�nh׾�#+\X���l�l��}��r�3}�N�:���sN����܍/���sh�fvUE�k@{(�
�y{e#q��9(Y�7~`��e�ⓐȃ>���1royt|��KGDD�&'��a��w�?�1��u��vT@CC��3x^J�G�(�єOC�_O�M�����^O�9��P�"��(Φ,��7�>m1�&�T�2�H�-1���R�K����D�z��z�;�����ֿ�^��#q3�S�,nC��(:���Ë�`��B.���F�o���Q*y+�0���~%U��)))HX'��1�2Vlc�j�}X ������x%{��ܢttg��ӄ�W�]�.a:
�C�<.)���ǳ9���o��}�~\�;���{���U�)�or�O±��z'���Z-A�Ji֛ݨ�-)`V_>�L�qy�ĥB11��$�����E�q�`��a��QE�	������xx�u|����꺀9�����}��o�V$��a���u5����e=O`���	�^�oa�V��+�HY��,��p��%=�p��O2^�ޠԂ`Fs�ʸ �|d��2�bϟ�H��-q��e��*�?[u��ݡ��KSR1��"��� �?w�8Q��`q
N��0�d��9j���C�{��DFFF`��T����]w�u��n��rYI����wж�� �&��f
9���~-U�������Mj����D����̙MF��}2F��1���z)��ܻ'3Kn�t`<'����f�]�@�Ysu�DH�}3�b2����O��/_�̸��{^ߐ�0��:�Dx;	��ݕtOI]}�����Ų���/�{C�V����m
����}���i�-b�q�^5~ZnS��Û0�:���ӝZY�&K VԒ�����@��b�w��S.�6�~��ш>UW��x� }�@X.�H����u���t�S�H��b��z�7��ha41";:�����"	k��<:� h	�oj4��"&F���`��0}ą,9n>MZ�/�=�ߺ%���,�	� ڣ��V���O���&�1�(~s����)��m?���R���X߸{�g?���������ނv�H\�>� }A�D���iP��6�Yמ�uX"��[muz�pE86�F����
(?���`b�BLxq~�28��o���:ܼ.�)$���۰���n�ET|O��mŻ.jh��y3,�[o�V��N�J��x.��X��a�x$���y����a��ک��F8�,3 8��zkvnQ���SjbJm!�+=CB	����|�ԇ����@qc�t�+Q3hf���V��Xؓ�����!ܴ%��y��r�������Ջ��sݶ ��&U_��"����������t��q��%�k��d'N㞱7e)�Y&���_t����t���X�7�LN*>����� u� �U�~��$K(<S�c��[�@ x� (�nU��&4�&L��4q��5{[g�����G�SI�1<�Jʸ��T8<<<W;=7W9�~Ǵ=����ݿ��N�06Q�E>���&��ѝ�`�=� _p4j�I�7���瘘��Ƒ�q�M��B�&��¶ߏ�V��;h�~K9�W�,�Ķ��N��BhȿdL�tk��$�X�%������P.[���B�>u?�o{�/*u�0��R�+���+~�jOA,��	�5�0������򚱩�Q��
������0%m�߷�V��)u(7E�S�W� 	��$�rq#�f6�cꋯ-R��mG?�Wz� >9O[���6q�A�s;R_q��CѠU��2��Kė-�-�G�m���R����6�,��0m���z���*�j>��nl �,�@�:�����D���deeĆHqR�2�Eީ�gbbHcgYXBfv���\{�~��3��1�ʧ$V��H���9j���!�+|������v��G'������bᐄ��|U��u��Qc|ͅ��>�(M��=<?�C�tG��!���_QۛI��ԏ�L�k����Z7����Rl��*XAz�r*))�.�|���2�3��.ls
s�N4������6g�f�c}�P\��F���G�1�o�����/��<�|!)���3��� r����佤�G�8|�!9��'��$&j��qdqN��rX8<V+�Bʀ��q�#	���v!���H��&���϶��LO�C�U�Ԙ�4�wu7�����Y��	��S����]�/l��ߖ%�$���-�.�Z���ub�W6��9�; ����d���p��uG4�z�Y��T�8�]���hۘ�����I���xxnx�_�Z�5.�o̎��5��J?�(4b�Y�4�Og�����=�"��_�g�G��}k�bYNNNץ�E��_����r��f���±uR%J4�h�<L3*
j(
E���M<�k3�����>�{�	-Y!؝wz���f�M�����j�%^�<��j���I�oe���o�K�vxԶ��(�,K@C�ihhڳ[��n�e	��'��#��m��qP��/�@?�JA��u^P�(����<_�KWRSKP;.�!�#�潎%Nod�;J���a�%s[Cπ����Ų��<���l��P��A�oA�hR1>.��>�{a���9�Ϙ�7Ȥ�OE�0�2��蠩�#HyZ�).Ge�f���W���<Ze���c�L�~9��x����nj߰�G J���TY�?��ͷ�?�EX��c��0�q��*-���"����kC����/�:��D�B�7Q�u� �"L��ʦ�R�<����:�k��躒ٙ�'Km���?����g͇q�a-�F���?}^C����9K����ab�'o���Ĺ1 �k84�̩MnW�Y�-d����f��֔ɨ޻�����f����+}�-�d�?~D�4kV�}W�7�,��9��j���S�0N7X�t�+��;9�5L�<8���$A���u�����ҙ�SF�t�A�x�����:u%��-��&wȡE�$T3�H���-T��6�as&�=��� �[�[�>n��,ȣ'�nm���X�p}�k���Z�b���ТSv�bK� �5��S{�|`�P�e<�^d����w�0A�/
$�m`г�����#Ҹ��4ג��`"&H�|���g&��YZ����JTn�g̫�i��X��2i���(졜ު	�i�ml/A� N<b�x�p�I+c�bB6F�UB�,9`������E��M�m||�VXؘAscCc� �]`���9� #��ѧ�����6+uڊ'��|���W^������%g�]41�q�q䡲�}$�H��:i�9�yG}`��2T�=z�So��?�}��qJ�6�L	�*kJ�p�[y�&Z�q
�d�UZ��r�J��(	���hR����$�ޞG7!'葏T�W4�Lm����E�U�g&�pX�V\��X��� ��Zi��3H*bQ������8b�v��0^��;�je0Pj�Eo{�kc�N�q�4>�I�K�y�>?y𦝰��笿�V��N2����<gc3������]Bs]Y2�(�MD�~DƧg�+#E�Hx�A�;�g��uXn7�st���.�� wqJ��]����R�1Ӳ1ǌ/:p��߶Q��n����v��B�"��y�j��x<�ʥ<�{�t|*	�5�g-֡T��{�g7����yF��C������_N��ҐZ���7r��&�Q��Z�t����z���	�d>|X��5I(V��bI�$q��~B��y��\^���Bb��z�n(��)̇ZF����}�I���>	�'��hC~�lA�i���Dw�1���WUŖ:����Z�4���h�M)�w�J93�2�!O\�'u�]Ƶ�{5z;�#��2=� �w���8SipS�]$��p8���ӧ����0"[�Z��s@�X�Qܩ��gv�~t�Q����1%����a]:��V�hZ���H�W��gv,�*�"&�F(tH&�)��ҼܝH�6k�$H���1��%ht���^b'�ثX �6#���=���ܷZɺ�2U�����z�pe&i1��S�Ŭ��"Urb�v�ٙi
�Ew��9�A� .�ؤ�P��܋��1r��Dh�N$�|�H��:
���=������� �j�/��Ic{00l'<��0���D�8�q��ﮬ�v�:��I�I�ɻZ�Ab\Lˊi���i�G�p���<)�oę?�Ԛ-�Lt��J����AM,D��}�j�"84����~k,���p�|3,�Ml�"|@����}"2��� /��IH����je�=�;�' X�l�V��3�Sr��H^���=H4�m����S�8�,mx�~ t
.b��g^��	Z��s�hth�¬�p�c��B��������4�v�ʮ��<��gl8�?�a��}O�|��j��K�MAx-���@�Ϟeְ6
�E}���6�\���]Dһ��N��|�#K��u�?�H3��?��G�<B��e���R����*N�B�b)�E���I9�x[jH�,������'E9�Gl��1|"�q�zI��o���F�&�ȟ<͏�ؿ���۫�� >4f}�� ����ײA�M��/f��~�Ԣ+)��?z(��K��ZZsb��C�C��諓��]M����|.^���.�e�s�x�~�/��� I����F�"��?�*%ǉf �Qi�+s�`EΜ�w2ӂ{>���9�Ւ�&��C
��-�Q9��*_����]`_�{!s�5����ك�0|4U���T���N�5�Z��ftaf���V�K�p �@�ĉ�U#�)�ںM�`���r�{2#�Աhnf�=�K$70�������A�ժiu�Z>G��W��'�������F�%+���������J�eJ��{�0��yH��(7^ML�W�ePh�'7H�q63��pM*l\b�/����V����/f������*�� ��t�u�����Me����8�ړ�\v]�^�-�zc�͇A9�,�D�����9y<'@��V��7ExPO �}�~���4���Z����	p��Eq'������7����S�[KAg�,5���^3�gn+��_<X�Y��#z�0$a�p�a�����e^XX���@ �^��i�T�g>�"i_mA�����ģ�~fc���/���JZp�j`�������Ц��=R�.g��ۻ�!�ܸ���-��,32����E���� �=2�<D�!T(&CI��4�[�1	fsC��yv���û���[~�f	�5i��DQ�ښ�;a=|7o^;?=\&y��̻�Ăd<uGGi�l+%�ĳ IXFi�4B���x�RW
�u7�����}fD�7�Y�F������	�棔R�W��׭4���e�)>&�<���aG9G y�`Q�ƖQ�H;���B�"��ZQۓç�,OR�־�SB.Hy�8Y��t�U�#�[��a���NO�|��}�/WW�����o�������'2uFdAM�3��S{�/i��&&'q.��Tlmo�����n\M��J�Zu��;�B6�u�^��;H
Du��s�S⑽�$@MU5�ZrF�(	���l�<��� ����}e�/��T���m�F�x��e���3�h��칬��xhFT�e`u�Q�Rx������3�m4==j���7[�	l�G� ò5��8oϔJ+[��|�����<�2> �]]���D)�!ss�SE�2�E߾�;���V8:9i��%����><T41a!ƽ��/4�������sR;���Nm�N���߁�a�;����$�c�����Z���~��=0܄ǡ���rN*����U1}Ђ�� ��Bj�i:<��HR�O�M#��ъ9F�ddF��`3���V����{59ƧD��=�����7uw���#�b������53|�T�ם~]y�/�6�K�2.u���=�E�����9���|�Eޤ��B �zd�G���4}d��x����]��#'**�O��G�T��� ����yO�X�5ɯ_��K��u��`�J�OD`��iFF΀A��.��6�o:,]ԝ�F�ZT_qCV_��:�U=f�ɞo=�;̈́zf�)T���k�+��Q��4�Խ����&���w���I��}y83�_)G0/��Me��q��8��uͭ��`����Z�*�������X�7i�鮿~#3=�j��J���8�F�<�yڪ�LG����%��<3_��H;5���F��h
����h6g�:&�����`�ZZA�^&��$)8�Q���'�k2d���}Efn.~��F���Ν���Pf��7�����c�q�Yɻ��]���O��A9�0V���+~"m�=��JeS�2䃔���ʵ��7�4�	T��F�)9P�����`! %CN�`����8$�����9��u?A�������5����1�tD:��8.���k����Ɨ��۾�����y=�)�f��:TЈ]��}��
�`�,�N��~���N��cL�y��|[ɫ]�4I�ݥ���'��dc�/�g����k8ҹ�s?�yؼ�0��d,�XG���c��3�M��o��[�{DU��Ə�Y���/�]�h6�8rD=k��#%l�7x�D�}��Hm�gӸh��KUrR��eԡ��v��'�p���'1k[I��b�ج���:�20tI���ol͈"ox6\]B�0H+)5ŕ���
D����bXSn�{~�3_<>�j�ɡ��\U�,D$}q�������1CGǻ����u��] X1N�-+h>@�c�
�j�����Ī�St�l&?~:�z�=c⚌Å�m����y��Y%Ay�+_&��6~-c�b�����ϣ�����WX\���u�t�b�����pٟPy�.`	
����m���+{����s�`k(~Lh��Y&I�fJ��x (G�1�"�=���ذ�am�����c��S@�u�ٚ*�r���{}�Fw?e��/���?%fz%�q�{RÍ}�q\]]�n���ѕ�@��>KQ�yɉrJ��������yW9[+��ë�i�4zfp˭�����Y`�e�2��3��`��y�p�Hd@�AG�N���*�p¨!	~��.�J�wee�0��}ʗ�e��pzG���S(�bb`��@Ӗ�A)�76\�2VN����������y�z���Б8����ŕ���&C�L�t�-����\]����0�j+��4�}莵�u��N��T1ʵ�"�'O�#נ�+�kkk�	�-׻^��e��Q�8�?��U�j��:4��<Cy�lI?�ƻ��ƛa*A,"�-1ǚ$k~��~d߯FZ%Nu������K\�]��ԟ"��oq�o�!#���f����NK�E�3]��~"�E����b^:_��#F�z#.����y�~��wa����[a��U!!��J�K-zl���oݠ�/�:����f�P^U5�8����t�&��[�_�#��`��"Eĺj'd1n�d!C�̶|��c����3�Vx_��m�����"�M�PJ���k�y�*��!�;���`#�?�c	��O��~���ǀ�*�,-�̥s6g;x��ރ�����h�wa�g�Dx�����2��ҙ� �ŋ�$�1����Q ���R�U���++H������U�����K�)�����,B��s�+K�M"�H�j$4Is��j"�lk�)�@�dh�iz�w�2����I�|�ꥤ�ڗ:ҝ�����c��c`����(E	h�<��~�g�r>@g��rT�A5�'�y��^���~�L�I����<�%�\�ϗ0���R�57���
�`;ZP����c�1%�O*1�/Fy��A�@
ZpLKK[̉A*����zP���"��?vK�����[����G�h�;��H��+�-�����$o�8�����*$K�5�DC'Pa1�Ç�7P��%�	_{��&�r�g�ܷ0��/HV��!��:�~I�������r�������g�~��!a����5?����.�q�2ջ>�¨�V��D�����m�~����y�:�T�n�ޓ�U�Pנ	���G)��5S?g~AA����[O�][\\K� ���@Ǵ?C���/�Ǌ2"�q�oߚX�"����^��d>Jta�;�/#m�(�K��i� �Sw"������"`�O�����嚹�4��Z�_z#5���T�ZA��FW�l��U��������Ar�|�8���ct��~��e��gk�)��:�n���dA9� ��
?W�GG�sO�ٜs++E

�����mMAx;��ӳ۳-�Hm���S�����z��ŵ��;��W3:����9@��c����xk��r��������Ѹv�žZ�N�8Imsh�w��V�槃!��Χ�Ls{�(( ��7J�_m~t�������w:(��� �#7u%񀢢�
��V�=��S�g�'u�����8���r'���˨��-���]�Ȩ.K����g\��;����A�Q�V�;���ώw��~�B��������VQȤ�)��;b������.Y��㧇� �O_2�ޏ��ZlfHV.J�OŒ���~3��ƚ,�$���Q�#JXo���
��۴���/9���4i�,�Lf@���b닔���	��l�6��l�|�4E�k�EFF>4���.��o�ݼ,P����AZ@"u�r�7��VR=�ӀN��c31�쳮���%���y� Ɔ��VVQ)1i�Z���w�1���R��N���s�� zZf���x뫾��+L�K���\��c^�7�&��aL�4
�$ο,W��]m���x�Xx��-�B��x�@�uǯ���7��]����_{d��Ccy�W�U>�:��72�ԯ�B��!^�TO���j���9��8��@gd=&!�y���t!p��~W���q�З.�"j���W8���+}��S[a��_��.v&��x�^�k��=As	

*-�>I�_c�5>�9Y�P&����{������4,4U5���)6&��A6>Z�$�|��X��e$R�u$�;�m*�2��	ȟO����o��3M)����v���2�y��.��0<��K��L R8[7�s�w=�P�ZZB�&�� x��Z�ȺZ�Z���zx^��>�zw�ek��q��+�䘔�|��w|���85'�PR���W��������5�?X%ٜ���y�����*��>�"��٫���XuY��Ae�"*fd��6��\k9O6b�?m���!rW��#Ğŕ��o��_�R��ն�UR4j�g��{(�����88��b����>S��9��G��׽�Fڻ��|���߶�e����� �2U�ϵ9��[W	a��JD	������h�Pn^ޫ����Qs�yyy����!��!5���H-T��폽*���_|��������MWW1���!
��<�ƣq�Ν�g�`�Z��1M%�Ji�${���T|r��j��9��Id�땃�C�&�a��Tk�􁴴�2 �}�.�it�n~�����J�C�@��	T�����8h�l��I[֩�ڧ &	E�7�����	� �NGۦЁ
	�߁�rg"��dM�C�Y�|bb	ΕC��Ɓ��:�z3���L~w2�࢞���GЅ<�00ں�ad�-xު����z�B����<�]3
����=nh{����w�5��������$~�4�����[k�#"���M�Dt�ӡ"� ���Z��*m��_C��8����-���+�g��+4��1i��rt��K7�q3=��X����m_av~����{ݭك�I�S���8��;���Mk��f���m��by��^�������~����Q�'��i�4���h3T�Ԕ+�[\U�gY�7=�M�lo��������4i[ND���`��z�Ff:�:����K��8�3I5�W�}�Kt��~�^�{�OZ�
s5ş���U�$Q|�`��(�~�ao����n������4r��&|>�n���7�QhXS�o�}�!88��N7(�}V�^Ó���|��
lh��.!A�= 6�迗���]�{��Z�)sL7�$��\�62������������Y�U�S����Y��+-S֩	�i����A�g|S�/�z��ê�\��w#��1���m�H�u$&:���E&��S��뿄��Ctq�-�ۄqW�Κʴ�[S��)_��'#@�-��Dy�W�[	`�<��Y���:j��������?��(�DXu4t>M�ʿz�:Q5�����Y>��� `��0Z�����0�Q� ��(�����-0�	�X(G��H̪�Q^iGL$$���Pk��B^��:؎�Pc�y|XY�$i�~?|��}��K&��ۢ�v����=������hk�C���tb/wX��v��E�K8E�=|vvFNْ3Bd8�\�
<�(0l'ܨ�}����`H�]�;KʧN1�&��.
!��<T�y�{��P� �h��|?4�j�����h����#�U�l'�ǉ��$v�f><1����P��.,X_�Z�����"�]��jq��/�:�0|)/�i1}���6��'�c�M�@	3$W#%�,�[�|�WN%�M[���K_�	��W>v�ѿ�ee�'�da*՝i��v�gD0�����*9}b�����K͒	��nsh��lG�:wux4@/�;_#A��B�V/\�]�h�~�{��v��t�u�|�5GK��/��g#bG�������Oi��XP�D��}���lh*6��y��׽:G�J+�ʥ����P�|X�~�9�X�����fm���#I_��*��m���999A����s��R��P/��+�.eTN�W�+ڧ�;�ƺo�L�#E.�t��{AR�,�þ蟄.ܵۺ;��"�D����Z���V���JK�J�a����`���C��β#���a�.�;5��&���{����@�Q��s�ďꌽ#V dpo���ԩ ���x��Wc��"h���}�I�|��������n�3������A�����Uϟ���<�ĜB�������_��Ӽ�,&v�%�UZ���)��*so>3�$���U�eP�`�`o���9E`������F�ۖ������G`����p��" ��|�~=��_��
�DBo�PY"�,f��0�N��tCq޴�$�e�gD-�����?����q��J����?dV#�X�9��ߠ{�(�����ⓑ%�X��Ru��I4�m�8_e~���Xp�Ǖ-�(�{��(�	�|�tg,(}�'�jH��p���z��O�S@���z|c���1KH�%ũ���aa�J�y�2���}�b�(�Sf��H��������� ��n��TˋM���W��Yc����|���ry��S��Q���_�@[�3�]�>�b͈_]��qT�
y�ܯ6�z�h.��V�.��=<R���U�B2��o߾��=DMM�W����S�$4Ĩ�|Sf32w�dǀyh�ó��G�LrΜ1X���2�Y��Y��~
��<@-��oZ �SqeuwCȰyߥA4��EfƷ��)-��7��IE�Dr����r��p�S;7�ӥޣ�=Օ~�k�u��������C��HO̭FJ�ۃ?�!#�q�<��0��v�	B��!F���Z,��.ǥ�F�q��XL[.�pjȽ��3��Wc��u��.���g�� ���hllm|{٩MQ����?o%�֭8gy�����-h�U�ͽr� ���c8pz�S�����KK˙ GkS��wj�h�-�1�笡Q�ѥ	�w��Z9�����!*H�L�_7l� �|Q����q��%���'WR�`�-����=ci�4j��V&&j��N�f�ȡ�V�*��Ӽ��y��4����m}k?�k����fH�
�r��͂#�7�kCy�H�F�������t2eeez��U�"s>V�"�����(�)*�@�Q���[F�i��fB��B��Ӻ�J\;W�eת���GV�j�>8m*��~#K�A���>C4��J��SA��]v��g�<&T`����@4�����H�x+J52�ii����o\	wh����N�κ�'�a�S\�R�uOu
Q[�E���U�U�:�n�a�2��|�8�:��?�t��D����Ƣ2����,*���Ɔ�Є�̘\�v��VX�H��d��m�`����^���e^z�Ե�p�j/H��ǪY�m`j{9���jYY��G�W"��޿���-Z��5f� �0��Td��; ��;�Ξv|��&I/��b���㣳�����T���Y��=�qߤ紁*	Jf	��8Τ��儘{ҷ`���l��>o(�o`do�>5��j�M�{��K<AH��������2�ӧ8�>�*hR]��a�������	��Z�������.113+����1�eI333�
�����C\��ݟ�	)((��1`��A���j����q���
�T�<��Pd�mߞ4�+�6�x���г�ӗ��7/N-��Ð��P9߯�f������5�㇞H��OP�����5�b�c<��]Jr0.=�E��mYt��,W����)+7^�� �#oz�@th�
A���Xo�(�2�N|�U�  ��$x�懡Эɰk]I�1Rנ�����(�d]_�����;�5X�14�[\� ��S@��pK�յ�����B�0I�U8���`�u����~{{�?#��yb���KШ����ݹ���*�����T��ڍ�e��)�N���hmm���Ȉ�!sۚ"����z�$t��2�}W_}�� =��_o�"V��ĺ�]X}��%kB�Eæi)x���f
Yq�H�g�h�ּw'�*�V:�����W|����߭��:���(�U�:c��ܴ�l%�@��O%�7�H��l�s�Tc�/��Yg��g�Z���炌L�] Ș(a�%8�4���<[�� �H����n/ǘ~9������������ܜ��X����ˇ-��7B�df�'r+����L2�e�����_Ŝ� �"!������~�@-��>�1���ɐ�����������uMgaiI��{r���5�w@�0�C��uS������?~<3?���3tk�0�����+Jʘ��R0������Xu�BO������TV�S��	�f��P����5}?�m
��QuUֶ�р		;�	�O�=��:�[D��+�탶��<���|�Ǵl���Ry =�C���^��3m�:G��$��@Y���Rk
�6&|Ym�4�j����P.#��i��jO�����K\$�N17z+��;)����T�ޅ��Z~�K���ᣔ:l##�=%�y���@N�Q��/��|O��y�6�(^�,n��APX߽{��ty�N�eY�s�ã���Ƥ{f��Ʉd1�C�F�`��1|��XO�>��ݵ,�!e��R�w����<pHOvO��l��]��[�@>$v���������-L�u��կ������f�M�/O�R��0� �T�@LD^vDS��K�a�m�od�F�t����4?Zz$�m�U�8�0����G�U�ׯjy�s�L�j1�k֍�o��G���q#4Oʖ'����G�E�=��p�2H���-?���Z�L�~�ז>���̳";(\��O���"��L�^hi��0�xˑ���
&�I�% ��*��T�/��Ķؤ$�ɨ�����iy���-��A���3���?~�7n� �>�1H�LH����K��_Dn���2��k��TpUTnе6��}�M6OS@SYsJ�_;��|�E�^{>���͆�����E*5N^�t �wwX��p�3hS�Q��9 �/��n?6�҅Ylv��N�5�G�uW>Ҋ���B+��[�����|�9I�);�r�-bq�5w�T���_{�Q�����;�&έU5�����x{@�f�Οvly�T��S��ĻE몕!�b�j#�D ��'f��TLL�����(��2Z�TQVT? Q�['�[�^_�	����s^P
~�:�����*����-@�,��:��I�RC��c�+��캶AJ�.	i�.鮡T@D�)Ii%�a��R��;���A���?7O|�����d-\é}���u�s�3D.)�t�ʷ����5;�(I���OF��z��%�������<��s��b�HƙR��W�o��1���9��'��8���P�F�&&���`7�M���h��Y��j��F����衖︍&�/���ǥ�����y�x�-g�Ҋ�ޓ�FF?������0~��0:���D'�]����@w�uLs�!��z4P�Z�tm����5ϧ@�����;C����?s���
�3[ZZ*�T�����=2ؖ��Ҋ@���*�-MT���ݣ�������-M���d�r�p��|�%>�^�u:]>�t�FKs�,zW���	7�h�l,B��;�8�9'���PC���1�3o�,C����󽎀fT�c�ЩO7��Չ�a�΂���i��!�|ɰSu����9��v�o��q9��U?�Ed�D����cX�ϳ��X��#���ȯ2|j�{�VI`���f�z���R�F��"<h�>���lEz�g��ذRRR�F$�wO�q?�l�~)-���Qu\�:��P��3^�����m�����4����ZO?@�݅o(%�Ջ3��\"h��H��~�괫p�����ZM�X}%��/��\x� &-w��S��){rM�W�1����������Z������sx^�D����u�v�?!�v�!�W����p �w4�cA���~���h9ٝ8��ԃ�����q�[�i*m�͆�����:�xӫ�7�u�����G}Q�{��c��O����Ĉ�Ӄ⃂���w��Ξ6p+��+m��՛B���O���z�J\�6M�G
4��X���kn���"S�&1�9H����?عI�ft�0���Ɔ#`5��dJ��r�����Z)	����3/���������44H�h߰j���Q�|�7޳�Ҽ.���k�n��������ۭm�3"��v���_�a�/r�ѷ����<b�H.h�N�2��DUͷ9�B����@87�I:a���d�b�>2�}:q8s�Ւg�_[���RI3{� �f�sI2OzĦϺ��	3[-qw6=I�T�`@@SU�#��NdoH���G��9�n���{̝�0Xc>9�T�4xcqpn��||�܆�zv����	=��[Њ,��;�� ..���
^��TQE�7((�J[q�?��!������o�IF����Q��mYߠ[�����'2�������OJMݵ��{��5m�{���|<i���t�9��_������i�H��$;{$9aюl%��v>����"��}�	O����f�g�߮q�X�k۶��ck�'O��w{$�2ǭ$��}[G����ڥin&���x\�~��I�t��9�`<��כ9����#Tt剴�l>�,j��9=����Iӯ���1��sf�M֫�4�6��{:�o�5���9·�rs�����o��zE��AA�(��]v��3/��sto}������x9֛�@8VN{�l�R���6}�3����a7Q�����WOܵ�ʺiT8��l�v���ʟ	��̓���8ը�Q�_��J"�INƕ��!.�G����]�+�y��o�}����b�(-g�������g#m?�dv��AfG�je�a��������c�Vt:��ʮ�CݘN1��5s�n}��2{�|���;�眮h����ͦ�� ,�Dߘ���ҍ��o�گ��dVX�ڛ�.�ѷ��d�@[����v�Z�nfaR������4�S�99evc�}��l��-��rrOܯ�ű��H�??jeeu�A'��4P0]�̕	�T5i�kWv���&��Yt�ft�0N���w|���&��
�P7��T���yO�u�F@<$���������4�K�C��6m t����)���{��'��ħ�qBc��빯��G���f�4&+�.JL�PZ�ܽw����=+���A�uoѮuӁ����i^nN�����B���0s�-�ev�(\��X���t􉾁l��T���9��a��7�]S��׷�2��FϽ�v�Z����\��C�B�	����uY��=��k��/�^��J�Q#ф��g�^�L�4��]0U�۱�Ap���)�]��*�����*O����n(k�:�E/G�K�1�v�ew�!�����u�-��˙��
�����8����dH�GW0���|F�χ�����QU���f�;e?�b�9����"��z89�^�kt���\�y'�Ī��aa��Z�pۨ���ZxD0���& M���?���8�Ag�;ts��rqc^�8}�v�����?3O3f�]~CM�IЄ̈��/�=�8��{l�!0Y��EJ�x��r��	=4�73=i��G����B��;��Ѵe����C�}<����޻��t?l��PSu"��n����V1$�S)k���=���G���{����hs�>�0�χ��2{�o��w2���6a�|5��Ľ�(��{�SqH��H� �%����U��~ɔg����:>9)��x�BRw7>���x��X�VʃxvL**����Qk+����`ʽݞ���~j�s<�Y��]\i��dOiA9��[�c�b��fsy��׭���fL�%�C�]mY�q�m��Q��k;�-(>�����ɈSɨ�5��n��(��ʶ,Z��ڽQ\���/�	[���߲pcj� �(�h�?B��)(�����20#41W�E�K���B��py,��6.���P�t�H�=v|�M�sM�P���T�D8c���1�7�Ǝ<�T�Rr��`�Y\�	$��q ��	���}�Ŕ���y��Sĉ�w�8=�%��[��gL{�o��'�����&��!����̇.|���8�c������H�����4�{�\]]��yQ��J�z����--O�?�5= :�sq;�^ҳ������?2]�Ԍ�C�UV�����J:u҃�ڦ}�6��� ��+W�U���m^���y.�=��=����H*��6p,R��Y �У��Iߴ\��Jj%���v��/П�&GZl�U _�|���S�c�C�ӕ����O7����q�tE�1��
*a�O��c��<؈X"�+ҳ*��J���I�ɴn���m���Ht����(��'�N��Y*�0�5������>�C���B8N�E���@�~[�§ ��RPP@��l����	bV�ٲ�9�=���"�1��^�L0��q
�F��^b��:�(j,&�ԛD���R�A��l9��퍤{�F������`yY/���Ni��(nMU�Y:��5L
���w8��(5_�j~w�q���h��p�6D�8�a+�&q;cH���)�3�� ���Ha+�����K��Ԏ�P4?Vг\	��Rw����%k=gs^Tkb��ϥ��^� x�Qf�Ǳ���FæWB�������q:��V��i0��qԬ�F��)(���\!0-"&����J�����:	�Xw���y���}�c%_�� ����M����)ǰ�eN9]׎L��+�V�~F�0��,���W��~G�|[��ɗ�r��G��1N07x'\r�:��1���-q�YCS ������.B�ӷS ��B�ÞEsݢݮ,UV[V$�L5���F­�(�5��R�.A_ `�9S�v9v�WZ��,*G�} �28�zh�L�����}7���4�x�c���5뼽��b���W(����
q@���� �(�T3ߺ8t�����O�doZ �C%���HA�#�B�vVx���ٍ�F�=��RI|F��wnJYM�<�.ծ�N 3�䓲0���miad�>��b^���^��g��<R�'�z�¡I�}!�'���B񎾿L���?��D�.Ui�yٖ���w�Q�|����aVZM�C�k��3����6?@`}�c�ӯ��4�3Jx�:�|����߭�%��j�K������lp��G��޳Ñ�ΰ��X:<��&"P�E��6�`�x��̚�֥ͪ��p�pޫ����;�sʟ?����E��nZ��&"9)���s�V:ך��gR�V� ����SD�u����2و�(3�IǳJ��u3+;�x�S��ϟ,���Kr@����z�_�Ƃ32A~FhѾ�qT��ф���w�Tю�������:N����"s����}�.#�.G�X�SI��hA�$�3���-� ԃ�k���r٠o��cA�-�9����tv�LY�,�Zv-�}��4to�b�ܐ�����Y+��e-߀A�̩D8�����O�ωOQ5Ǖe���%��!���U�E!w~�1 �u:0��%���`A�wO��Y>��u��O�OW>(�(K5�/�/z�N��!Be�|�t��h,���:3�}��f뇎�5�8^G
f{{6n��� �-,�b�� ���g����Z��/^��D� �K��Ug��T���j���CL�H��c��m�~��T��;�S�5M �x�K�E��[�3GWI�����3�oi�]k�����(��K�)��}�+�}Uo��ܽ)0IX�Ǡ�q|w&{/֋���G����c�ښ=��&V�0�)��m��0tά��ߣo�>�A$(A�T$
�Cы����x��M4������$���]�:^��̈́)=�*Bf���2�	���� hv�?�2X(����)�|��_Wz�=����cI	5R��
��0@�w���]a��<���=�<H�a��s��zo�۲м���+��NL? ���n^��]�	�Bk�� ��c�~���gG�H��F-K��p��Zم:����N<q�/@sNŜ,��Zf��z>���?��KY��ڷc�}�6=}�$�F&�d+��V1���,����U5a��I�����B�/5�0�*2��������uc�U�{�[e�^Ă�}5�e�|�L��FN_��2&XlF�t��u������>���*�}�'@�Gٲ	+�9Y�]%nȓ2(�>���؈|n��pp��Ѹٱy\�̌���x�D.
!l=��mk��]��Gj䢲���L�('/y�����y;��	Q\*6��M���t[ �O�t�z3$C��H�d�p���_!��ll�6��I1V-$"���s���0��e׋r���%��0�z�ذ�G��-x(@	�W�αJ^��O���n
lF��n`�<.�E $�^���-l�]���y6��[}d2ez�j2}�\�\�s�
Ec���;����W�4%��_����b��&���G?�k45'�j^��D�����g���V���R���ϗ!u��/���.a�,�WM8��.�	[�0	^��R�>je��z��T���I���bqq1���|����:)�%h�.����xz����ެ�P�:R#����]]��Xd8l����i[X��jZ����FRYl ����H���qh��s�4�ʡxb��xba���u�;J��Ⱦ�m��G�_!�"]qc�KN��E��{#1���#E�o(�.�n��3����yY����%�R�)"fV��۟S|��>��Қk�^<�R����υ܌\=��X�K���$��(���ˌ]�F���|j��Sb?��ݎ�أl=��Μ�o��5ۑ�fEJ�9������ܲ&��4 �� ��llHAȃ���Ζ7K|���nei	x�cKKv��%���8�{j�]���Ҍ`�i����I$�?��t1�V���>���T�6_��ݜ�����۳�k.��0� ��ƭ�	���Q�������|�z�[�cE.��Є}5U{��N���)�!�~}:�����nq\R]#�����e��S)������a����-1���p�y�
a�R�r���;,��|U3l r�9���*�O�Ý�~ݛnb�Iz���z���e/�sz��%�-���j6,�w�u���!ֆ��fE���"��A���`:����',��!�εX��*y���7}�<vE��S���8L@5�Ʃ�9�����%˞p�4�,;z�y�8�v��t��
�����H��֦����x"�Ŀ�Z��%/�����ss:��l�v��_ۚ��a��d�����e*DƸUJ�W7���.������[�����P���˫nپ����ܳZl I�~��-�ϲ���~�Y9��3Hs���	��'i�����;4�ӻ�2�ڄ<z��{bZTpii�u�&�b�\� ����kՀ2�S%�����E3��%�А �NAA���Mߊu�#���%w�0k@�>���p���Iq!f^į4�ù����]~�xu��ub�@|��k�E�W�hÿ�Fv�җ]8�uZ��?���4s(�.0�-X$��Vo�}�H�^Z-턘�����o�?e���;ψ�B�+2L%�6��{��|~�ӶMX ��S�6w��5I2+����L���5O��S�g���gt��9����>��r�Q���c�ҙz��?�X\���v/-N�Vʞ[K'q�,�R/|Q[}�[ɧ	UJ���Z~����66>���>�H����噰�A���u�����z*$u<g/�a����9U��ڶ�[��3��4�Kj��!�r$�e�� �de�I�3�~.�;ZCCVK��`ʖ`�4:`7��~^��Ҁ:�W��Խ����){�JR���S�������0�K�z�ėr
�+�p���Rp�8ѿ�ym���&���O�7�I��^�h�V�������&��}��?<��:<����8�Ժ=�����gwJ� ���[�^Vx�,�������?-	�,ŇZK���}�Qh:(Dc/���n��8"��5�;��5N0".�U�#?TWSyyy�l)BGu�A�S6���ԋj���-����/J>��W�PMP�w��4���
w����!�7!a��EL<;���]��O�G���M��D�-��dFOci�p#�7�t~'>-�3��iW����c�'��H�R���t���M�a��W┐�I� *���VU�q)l恚�V���/�:�N��y�S{R���}&��#90�E%����Ԉ_޵7e�.%&)ġ�R1����t\+�^&Y��Q����M����6�m��)e����CK�4�I:�~p5�Pt���w�æz��)���%����*�ҧ��d���1�k��u�c�{p�ڌ�H��&�׀�����*T��d�T��ƥRrI9)�а��S���a+'�P�C=��*�w���m��3��
ӡa~�.��}�H-H������������nSw��k��3,z�B�7��k�Vq��:�t�H4;m,��0���MJ����uy��O�q�H�����1kuX��x�70okt�,�ǧ���ʖ���ͥ<pVR?��~{��pw�(L����ăɲZ˝2޷��w'���T��9R�?*D-�ϰ��c����]"|g�A̭��I��Q�/�	d�A�:���ul.���\/�)y5v8;4�����_�\���;1d�C�m&�I٣��Q�F[�+����."�<����?�a�d�U���I塜ݱ�N�oR�s�O&]��%�E��j��k�(F3�M���mL?�O�^ܑm�u��:�b׌�}���k��R�%J <����KŴ5�,�Χ��HǞ���U�Ũk�򻛻��\����9پW`�E\�)�1�uNk-3~x���|�����	���0��}g`�-τfM�[��&�լ�F�-/���	���/��DE�o��WKlw�t����TU�E;>��a�NսC��Č����^a]�,�es[���:������5{�!۬�}��L4� �(���́��#;���ΌJ��'�B�ڭ��d�|�( >![�o���!��5M��ׅL�
3� P/z�bnA
$���I�p	wn	W��y��@9V�K�-�d��k�B'.55�QMkJ-ʙJ�L�uf�(�k5�A����)���ӭ�t���Ũ��h2d�'H���1�T
�^���)��3~(J@�22��`�h���������,��k��I6׽ﳙ;�%���z<�r��F��{r��P�#��7+m�>��$�|R6�܄D<k���bvO��e�Tt��2l{Ε_H����v?"�H������bg:ɣF����(wW<��]6����ZJ2^7�TzmZcbp���K�c^�y��1G�m�Wt�^�]�yߐx�J���/���h�����)��� �my�b���?c弡,i
.�@�����"�G�#I�e�:�y���A���r��!�����O�7$�#��H�L��������Ԑ�9���+�@TM�/��Ě
Gd��k�Vr,�w�%��V�Z���G�RH46kΖ�E>�=�V�i��+]���Ӂ�ܲp��_#_�M"$���*��T	+F,y��p�veoi��#BnY�h?.��!�K�g��i��QUs�SQs-�����l��T~�W�Q�|���u�,=���0}$A�m�52i{��5W�C3p2ᾢ{36_鏘����{~�L�;r#�DC�U+ӷS�K^ߐ��\��x2�����l}��+���G܇��"J��l�b��e�������<�|1��<�E��T�r�+/YM�Ƒ�
�kF�]��0@Μq�8u��K��Gܞs��E��S�	������5m��*ߓ z�����J~uv�7MD�7<�*�* �!RZh[�z}�$�}J{�N�G�����JĞ;ȏ�!��R�~� BQ�����=F���{D��]�:������L�i��鼛�Tq1[��#ED�L�;?{����^���v���<��onKS�FʥG̾UujO7z��Ҕ�l�v��x�'��=��io*:;�X�X ��w�%�)5_͗�������u�$\�-��[4�"�h�A�\8�r�����whep��ܷ@�T�������}1EM
�V;"�#_?)��K�������*�(��'D����r�#���u$�W�ݬ���xS{)����mv��w8L������H��cg�YGN���qG]g��	
H�uA���@>&$��N��
��uJ$e?c���p ȮO��+x�̈́ٸ���a�o�I��uӐQ<�j(���]����FGk��utJø߹I���J��!B��6���թq��(Uu?=>��y�Åm��)Q�jq�Io�ב���o'�#*r� ��3�W���qun���&�6�G�A"5�9?vҩ>�:��v�	Ju�yd2�����3h�юV�C9��t'��[��ʦ/������9MXˉ����=Bn��د�}�c��7hP(�e0`���#�� rs<�|@==:u~9��#[:$/u}�T���h��>)�H;���+&�Z�S5>\���u`��'�։������sxz<"z0�tJZ�fm7+���"��9,�̾��O���/�"�"� ��V���Yg����Y��]<-B	��I�w[m�����4�6eY�~����A�w���ԍۀ��=�v��p�����B�v���
��a�A�CE�P���V_9S��EB��E:�!�,���s�4�E�>] U��tD�2S`Aq�(@�W Ջ�P�|��%�|(�]�OW(_ݐ��+�z}����Ӻ	�8�v�����_���b�W�>���;F}����'I�:�?�VR~smO����>� 0���Ǔ�MI4�5��s�H�����q�0�]�J>+���~y�|��k��/���'Q�V|���R���߻���c�(#����A���j�ܐ`H�[�������鱌2�%Qΐ0v�|ޅ���	}�w�I:Dt̕�S�LǾw�%$
��E�e\g{@����ɦ�G�In�q3d�z�)�e�H��4���p�-֜�g�=�Ҍ��#,Ι}ݺԡp-��L	7"���ܱ�1��f�z��$�y�T���٥+�}O��aa��Ӆ��`H� �C�z<���ʅ�u���N�]�~WMf�l6�Y��[G��-�����Ƶ.�!��������di��^Ak�m��~�hf��:Yr6C������a�����_��c�a�@���C�B���2���F`_���{�~�4[�Lf:a0���Z(��d��fωMɸb�Y$A_9\Ti�4<��D7rN���MqIq9x6��z�9<��^�+�j>�:�R}H�^qb�(+�ݾ��O$����bO�s��^H ���tW�)�z���4�p� �?�:	����Bc�38?>^�Cpw+���j�þG�v��pH�qڨ�R��Q�3���n��8v�0���>�����_�ޅ��AVI�I�v3��W�:�A8��hWZ�z@�{�
̮��J�8��F�Z� 4��UywZ(b$�ާ��=�st�<��}m/\��o��xv�������>���#8�n�K�T�kY|tㇵ)�z�%-���;��W�畞�O~�#C�(o����Xl�Lc���;*@���_D�ʕ890���f%�� ��	��ٗ�ެW.Y�gƂ�������5�5ȯ�x�#����@���������y�׸8�A���6>y"�M���s�`j.��}U�<3db�0��T������$&y�/a����;y��E֓���r�K�Jf��aX���x���aJ��J1=���lc�l�Ӄ�s��+����άC��t�V�)��6��^������R�w�G�G5$��-��%�<{��L(ɚ:�1+٨��7Jn/�ۏ_�EO��Em�ʢ�6���>��9��(��pg���j~;���Q=�_|n���6�&�N��@P1�È���0v�lcT�Co zAL+GH��@{�X�B9�	�߾�vT�HV^��8�+y_	:T�e�b?����iP�Р\]LJ\�8���w��*E���w$ɗ2��&hMԔ�M����`���`Z	��j���տ%�.$Q�qW���̺��i���~�4ZˌK��m��W����B7�R��������<?<��X��֮Y,��z���DTl�2�|B�Q�h�P=�H�w|����7`� =�ܾ"HO���S���2|��~��ҷ�I�w@s��T�nNn��"����|wV'ȶxZPc�|����IpJ�B��0��~����Z����`׀h��7aJ�E���ޖ%�"_��!ucQ��d��L���pr��
`���Ԩ�0-.���%j-h��i��ʺ��k���WFo�L�LW5O�M҉m�/�3�T(��a�>��h�ف�Ehe��,a(0��z�携o�z��K���#�eP����o��S@PB�ʎ��)\%�>�		�(e��	�gKu�S�Tݧ��5x��(����7w�gYr�k7��`�$�-6��j4%7��M�ě��G�r�0���h�_�\��($$��*ʮ:��giǥP�L�S��=j����;ymk$�78�⟜�8	'���Et����<����zR���M�`�Ě��NŚ�D�z0��Q-�e���_#{���Ʋ����G޿�M Z�ޭ~ 5U��Xl$i�h��(v�ss)t�l4�N$����Ƀz�Y���3>��,j�n"�{��9ݝ'?�<PV�I�3��j5t�˔�����3��TLj3��;���T��b��������a4ߥ*�ޱW��fP�k��%��q�2x��?&%����
���u� t� k���\�Zx�iil�
rۈСh-@Y�>��B�O	����!A�����y�<$j�:���p��zV �}93��vH|�����$��_�t�[�� Uo��g�-O��T�ri {!���A^���9�D��C1�s�a�`'��*٠;�ldW��0M����,�}��Ǵ��+�p+y��O�,ioW�����fx@�I�}bt3���V����8l�W�eϠ�O��>n�Bt�@E�S?�fj��y�ة�+}Ι2��"�!4�囙��b�S���j�t�qj�y�I'QY�v�⮸�%S,��;P#X`���w|� F�tG��'��6w�륻�j�&R���ɚ Dp��
]�r�+Ԛ�p7;��̫�ꟕ�Dj�P���Ϧ��z|drd��A���=�O�p`���s��D}�^�=Qx<��A5_=R7t��qm|gI�s����d�$_S��B�S*%��B��>�k��g��~F�Հ�~&����`�H̋����v;�̴:��5��,"� @��pD�0� V��_X�#E��)8�h3�#�pW�P�2�X�^�p_ma���~b@�-�I��F�bA$���ֻ��/����7A?]ې��|���Qq@C��q��Z]������go�o�mV��䀹U+��9����q.��.$ CC&y����-pC�JU:��M�x��F��\��D �'+����!�s�K�6�l���l^n��2�<���^�_�I��d2D!�`��z{�&�z.ʊ������!��ˇ���]�c0�f3�s^*�N�B�qE����h�̊���	JǋtO����h��NeE�t��T������"IY��2�P"B�[�Ow��r�v��2�"�����??q���s?.1��M+yiڬ����uEz<Ж͐_�w\\ м�	622��ی�<��=~���hS�-&��V�H�T�ID|3�k���gO+^M�p�w� �tn2(M�7�H�c�9�A��1���Plb��b�q�!��w��j$�~o8~PXK1����C���my�`T�&Wြ�'kM2`h���Հ,��� ��\8�IT������X�z��u�H�[nK����I9�s����x�R�\��wX�㎱�]V̩�g�r�B�	����PK�#�^��YE+S�w)����JNtfTߨ0������i���a"zӆ~�9��QǝQ��� �7}��A��2%J(�c

b�N\�6��0@����6�����L�XlC�؁X�z)(*_:
Ln(u�v� y�.�r�l�I�
���_��� ��5�B�k�	������/��"IW��аTj8���B0u��&�Թ���^l����^v:��A��)�f�L:^���;�	�7�F,VO�x�*�u�ޕ/x?~���[��8���3tB)a�e:m>N��m,�$� ���&�q��U�� ��fv{�]2����lQ�KA�����^	�^��������F��<�G����\�z���WI��n�U+u:�ª,^:��ן�x�~�DI���� �3'�ȕbh����1��uV�ꫨ*2�.	X��K���tw��sZ
,
�X���W�y���H�Ǣ���&��"��n���x2�.�����M��a�����Ah��{Q&>�#���=a���q���Avᾄa��*����H��A�ֻ~�B���N1{.�	��"r�
D���vd4���N������v7���,��<�PmO\д.gI�]0�$c}C ����ɋy��yw)�H.nn�j�'��A���s.�tC�"]:k�r{���ӽ��F�	��֥���F+o�¬ÂE����9��� My���@Ǭ�3��\Yd/T���� �..#��u����}t��)&pP�x��[�[X	й���E�q�l@qaaK٩i�q)j�q�����irG1R��b}����Q�6R2)��+�
ʩ�/^�p��_����Ύ�����`�y9t�C��
Y�+@M�����v�J�vk2B� ��(K��/9�IX4�F��)��{�봈{�DH���P���8��)�}���"e�=������1�ӄ�"�/]����>d��{�E�{�-���!���7u��sm���c���]祐�Wq&pc"ҾD���Mͷ���UY�)E���0+�����p�&''g��a����GcC$e��%�x�����>c��Rc��@7<7��m�C����8)�E��R)F��^�M�i�֏(���4;M�U� s�%�8�`�;�F�D�a�ʵ�k�?�}�A���4��Z�p/B*��_D�J{��D��kӏ�䧛sm:+`p��1���e���
Ea=�4ȫo���V�W�Q� �2���ep����Lz�lt����P�U
�Cq���Jh�����ާS�m=������!�6j��Ar� �"3m�&��L�v�b.��Ez���Tu�:�����׹a�ʈ�:��(��I47��a�yi��ì��Q�Z|�G���Y
���kW�|�F�*�P�h�go{{��ox���i[�HD7n�W2��D)�b�
��rt� �G�M�Pa��[��wN�Bg�83����#WQ\����,�LM3є�����M��c�v�����|��6b �6�X�X[=�*g8z��Ά7����� �1���X""i[a�����4�J5��W�g����x@��+��f��aD:�}H��]={%j�J�$������;��2���ip��Hп�`M���}�x��Q��蟧��+͖�J�	��me@ ��:�.ht���	�9�	�.�.�Q��/�7�^uӚ�պ-�.����G�o�Z�Z���3&'i%�c�\��`J�&J�q�W6U��ɪ%����Թ���p���!m�� {��m�4&3��`:RQ�ǱV94l��m�r t�D�ldѸ�S��Su��i���?i�_�ZF[�׷�Ps3��}�
g&D�M��^��|z�f$���?QBW-��$y�~��%v_&���R÷*�`)[^!��{v��'�:!ۂ/0�0h�I��7'����M��ֲà8�������Z�xK�GvH��s�K\���.$g``P�ԤB
�$$P׍Zݽ{ȗ�1�NM�_��k�D��dv�x�����Fw���><T@r�w��
&P��霻CSR��d-��1��"yq���
D�kᎤ0~ݬ|%Lnh��7���dCk�3}�pj���z�����y��
)��8C�����&Į���E��~�yF��Õ`_������8ǫ���U������@��ih@�����;����}:.M�i}}=G���z>%:�q����ɱ������w��	{'���sg�9�=T���i=Q",H�Ю.����֖�piHa��!�����d�(-�+P�����I�xN�gW�F8/��X�zR��k�|Q##�+�A��"�J`#��_���#�׃D&�������[h<	�4˔7	>���������QB+;�v+.W2�F��Ϡ."""h���� �[.ήe�&%Q��<��PQ����w�.�]�}''��㿞h>7y�k4V����"��?����^)���G	-4Ao��䏲�^�WR�bna�b}E.����Q��R���~��)>)�Y>��c;� ���xw�#'".qy���y`Cؘlgo�:�����V4��A,��ob(�7#�À�\~���y�ɠ!Z|���)h[i=�����Y���W��?�|O���6�zc�p*��f��9���R�����o~�A�^����]�X\B�VRR�̰f�R�xH"�ul���S����V�y���M)�K���`��X�������H!��]��.��w�F���̀���޼�⎋OJA8=m:,&"t�&9쿟p�Hh�p��
��8���$0�h�5��#"X4��	�EEAC+�׿���'
�8S�%Z��8�`�Ä�����ݫБ��$Ѥ���˩������e�Z������~h�͗4qm�����3^�3{�V.���f��^��%�I��َ�t#>�Y|l��Ի�t���׭瓼�'��<K��L���Oњtx~덂��:!�/�������V^o�4K66c�d��~���-n�o����r�~�M'%%���߅�b��XF�1Ա��߅w�ͼ>Y��EWY߇QQQ�L�x�|�:n�����D[!����7�=��#B�`v]V���o��	T\׊k{�\�O�xpٚo����A�[���<8)�{�l�h�lG�w����P$��/c.���ZeM�mc�1��V|��ߒ�W<��d<���G3��F\��t��N6{lb�7��4����~��M>��LZ	�JO�_�-���^�͗��:>��k�0��If��%z8���I�?���@;�����4)�[TQq{�q��F���.MП?���_D2�J�s=��Ƥ�oa�{uXX#33'���G��TӪ�S��ϟ��\덧_�َ���7N\�Q322����Q�6���?�qC+�.��<[̀o��v��1��[���%ݞM�L��f�[#�����R���,r?�p|x��P�8�������n�	�7������K�����-�|E�=�up������6�6�|֍���M�s5EC�tG�>�LMa�Sp� X�pdl�����xO�z��'��˶���\��[|�x*�׹]���@���^��q�[9[Cc#�gNa��H�F��R�h\�H�l���դ.n������R{��]5ϧ��?�����4��@@Um��׸N4[<D�c��?��iV`��2Dz�4Sn�d�����~�0��ZȻ~�3�/)��=n�˶�'e!���9`;�ޕ,da�>Y-d�9�*?RLl�g����\�{w�|�
#��_ZЦ7�)&W-�,�������Ao�ͻ#�s@J���{���. ��UZk�����a�}���]�9��fg}��]a�o��9Q�� e?=^OO����@̣B=�L����v����2�)����%��+�q�Q��&\5��P&�|j����'[m.`�˾�M�f�'�֧j�2dR�	���$P����D[[P��7�ige0�U+	A��ׯ]�4=�3���lqi����������sv�嶶ʯs�q��D��}�c4�')Y����[HuCCC��,|q�)������릑��me7�����ǩK��ܙ�ii��=�)��s�� ����
�
K���@�WǻU+��@�A�|��>if�;N�<�����T~��^ȋ�y�I�Зe�W���⫝&�����Ew�Hƿ1�љA?�ߵ�s�y~�9�/�g�Ew8U������Vw&�n�v�l6����ߑr�$(}v����������[��n�x��� ���:U���nH���K���ե�y\��Sj-��l�t4�t��'��,����)��I�~/��������fY�M)���AFV�vz�=�&��N|G�`�o���=��l�>eȰz�����P�S3�3���s�O �T� Jɝ]M���&�X��X��<1���bO��_���z��M���c�+O���9�ק���T��ku�H�_i��\��bhh��qqn.[ƫ���M���c�v���|��j�'��F3�`�OMѯ�G�����W����V L[[{Rw>�� �s�~%��Zt��߿�?@<V�� ��E���;ou��w�nmBB�B��dm!e/���%ٳ���N��Qdٍe�2f��Ԍ}c���>S�u����9�9�y��9��\��z�_������md��h��:� �E��^ա����/.�!�!���3�A�ف8�p�:i����lomZ6ň�	X�������7-���)��$.�:v��9z���@���Md�|��dd2�趻AY$ '���#`Q�����H�HHL$Lg���(��7\���;UH@�_bs�) ��J�Y�o�~��D���K'e��9\����
�Z�������;�w-.�����/���^�k��u�Vb��C�%|���b���Ì�k�AN���JOp�l��t�Z y1�j6�
B5xR���a��F���&�-�NBB�A0%4<<�$S���"y������������Hf]U{{����J��׭{w9���R9�� ��!��5r�s�����)�q����\�
.�r())�V:uq1�Ʃz��+ܛ���i��'�՟���Bv��-�ZZ^���|v�]�����������?��Q�-�_� "����$��=`�IcQ���nH�ڞX�$O��`�Dr���@���+�Ỳ�mu�Z��� ݮ�i��AL�cQ���4�u��rJ��q�5(�߁9�
���xLmD�{uO�ٴ&�������o��Ehá9���eȌ�)m80$*i�ML&��(��;6��
���H/|ОZ?�j����$��!��<	(x�o4�{�'@�O=ĥ�V�{�p!��{����8�U�����J��e{��K�������@��K� ak�H�&j~/����o������n6�rO8U���J\�ʥ�H7K�* '����]	]XX�"ձZ��|]�[d�/_�<Uq��ѱ$�;;�?�MO0%���1,�HX@��+v���T�E� $����AX����NK�Z$+������C1���*$1GIZj?�`�-�7���IK��/_ު�r�JQV���w�[F��\�G�P�m����q���	��!���⎄�s������@�睙��&q4�����ÿ�{̨������ $f
}7׼j9F�@
�_�Mt��ý���'2��%���- �d��8ށ�Ds<3$smk�hjj�W��Vd^���J����Ar���,d )�6�D�,�^ɱx��� ���� 6���.P^,��������lI��lu������PB��~�H��k�pK?�W~G]kZa��xKH(̗�B�]�,��^@�7�~z�����ђ�Һ���u""�A���Z������7�^ѳ�2 ���Q$^�-��4^����柡�vn��K�}�	P�G�u���]����?�?Q��� �����?�i����=�:������Zɋ��T��M��}�}�ξ�u����+��8� Jκ���I�.�N���ځ����c�bΌu3�SJ�_���d!+a��������8��Ͱ��?6���'���mn^^X�m�ۿW��~�b"+��(��|�ĵ��z�۫r~T�?�"ۥݰ+ՠ�S��S��^	0�����X��xS'�"��r��߻��\H�Ǌv��w������7��5�>f�7�	�LX�OW���3���Ԝ/FWis}ȹ���B'{���<��ia�F���Aq.����s�Zp�v3v��d�p�^"����k�y�L�ut��I���V�(}�c?��IG�U�Km�;�ַ��_J�~� ��ȱG8�i�r]x43+�oS>++�G�7O�n�BD�]����#��M/Po��F]�<��`�P7i��!vk�1"+�޳q�dϫC<H،8f^ű��e�����M�Փ�z�,��4YX�U9'�]�6v8��Ү�r��ҜL�N�;�J;�_yyЭW+���%=����J8]�t�c^��x��>��_D�?ےrIǧV�3�r��@WS~M�&�D�V��F^��@���%o�G�f�p�(�6��o��>J��:�ٺ�mR��K���G�^���=:��#rS]u�B�fQW�O}l.�f6F�ȫ�*�{����]2��V�:W#s����9�H�.�1<IH�<����#����W����,V_��=2��[{�������nt��N���ȭ���t��C7r(Q� ]�Շ%&S"�h��K���2�%��P���M�	1Y���/��#l'bq#�<��eE&���c�V^no��*�190�aD�辰�o��	V�;�ؑ�)���!���|��1ޞ!9e�G��X�v�hIA�U�B�j�׃���]�q��Ѝ�8�2^���� Ka�ۡ�B��֑�ٙb����Ɓ��m��V��+�/P�f�,E�ڇS�){ߺ�%��#�g�t;A�0���~t&Qv#�\�2CQy+�6iv�����@{����|� �z���j��^{�3��88�)����a��iᤗ��*+�y���9ƶ��3Tu�Orw%��{��#��t�}�{�R%H�Nl�%\�Ԫɭ��Y�c���3rxY�X�ꊼ=
�G��$�����8a�HхK� c�;y#�11t�u�����#��pmS��D�{~^����G�m�������Ǆ0�!�Fn�d�-�m}|V�;��	�`~׽�#��{#Y�Դo�������>F��U���)���&񗌔KMw��f�����fFҝ:���C} �CyLS�6C+�&�.�Ӽ�).�1􆄵����KC�ڊ����n����]X�2 ;�K%V���8��U��O����T��`{��U�f~�V�zd�(|����s[n�A���RH��b�������o��Y��#�-�JA�"+�TVF����5vy�b�r�,F~��GW!W�J��cs8�bp�sM��7M��
&L���-�~ߴ����!-��ɢ|ٜ��'a|]l/��n^Ш��
>`�.g{x����
e0g�����LR��4�	^��&;��@Y'yw���������K�?�����!��]����t ��^��H�:hJ=���o����=v��7/��<���ЅF'c9?brqje��(��0s�ied�&6�{Oɍh�����HԾ��Z7i������9�,��OO��P�I\2��Q�m��B/7I�U��/�f���t�)n�P�'D2���ߖF>`жjY��Ab��!ޒ�hlҐ��wU�7r�����Ϭ萕�[��ަ�9"Q����I�7�Lc���������)��R�f��M����2Y+H��Ss,Q��,���
@��υVB���4s�<*-b�U�6��&�)�qlާ(힏!u٠s"�����vxh��Μ)kG7�1A�����T��,<��I��K��W?��a� �X���O�u�ǃ`=���^锔�p^E�둝i�δ��;�
.�q2�P ��=��7k�4���_���L��%%�婝O��W�\�i�|��U���hIY��<-���ڊ�����ɱ
ۅ)L���8F�'%h�����8[���\d�Cu�$l�
���/��0Y���i����D'(���?��ھye[���H��In�a.����$E���K��(Q�hk�4�5~,B��653b�^����XO�!frTVvDNp=@s��5��Mcg�+�������A.mP�N��s��Ϯ`��Л�|H$`����VS3E���ńJ���ۅ^N+�|�2�T��
Ё�!�}JJ��'w�6~�. vFxnp6AĲ����9KokV��q��T�S�c)޽(C��ut�+�tA��ܻv�P��ϱ�$0�2��xM���pz�VĨ����T)x!�X���,��; ���䢽}��#c󓼨��i
��0����D�%7�����,3�
��S%D�Oq~{v�.��.u�J��^{���R�ڹ�.������sAYHy�k�-:c"��}K��gU.�ɜ��p�0\��wmR�+�B��l���2�>�Z�.bP�}��9؆-L���T��qjn�J�]D^� ���%qfnlhHU�
� ;zI��`m�IW�qO����fk�.��J��r�τ�W9�YL�N 	��8�\���.7B��W��Fq�B�|5_W�^cr���q��ٱ�Y_�c�Y�:W�vt� �z'1N���ஃ6 ��m�(�!��(�\������+�k4Ϣ����5T+-��!�cTr�Ā
*Y,V7�A6�S,r��iJ�-S}C}+���
L;m;�GU��MVV�l�,m����%��&�I80j\�Y�Vx�(��G�@8#�_��">��d��Z]��v����Z>*#Y��Q7����%��$�e��/�'��{9�wj;Is�n�=�7�����U,�(���(~t�T�� $Q)�>Y<"�s��^$@���>lXN�Fe�iX�_��-&09������Ҵ�ŸCN/Ç>�5 >�� �V��zu�dS[Rxİ�h�+|R{m�x.H�d��B������<�=:*����ZkjY7xP�T`��Xl������c�Y�nV~q	C0���)��^��t��*%͒e1|<�T���an�}D���cB�� �mu�jb~C����xx��P�sp� ��G�����RW�[��{��ʄ�F	��X�vP�Fs�-��ѤT�|f����C��d7��U�V-�}��I��\!k�>��Q�0ny�.��O/��<5��抣�QE�ؼP��n�c�68��;�N�R�us�G���_�r��|{� p�Ip�a&tg�+�3��Y���a󾺯�s٪xU+��o����P$���u-� ��v�0bF�:g���s�[��PCFta�E~��1^�hA�1���ګ�qG��K<r�`*�g[��?�f7b)���r)��3yke<�M{Фf(`nmA.i�#w����Q�o��,�#(�hN]�\�2;� ;2�j*�U�aoXX�����D`�B9&�u�{��x���Ģ��>N�~^�xE�m/�k��g�4�'��v&�	��@�����~1��_�J�z��YbJ(���A#۔e\8Ne+�T�[l�\E�]���Pt�2�f+�_�Q�Y$�/10_��=хھU�b�|en��h��k�Ӗ1Uq3��W���k(���+���2zT�Z^����Q�i�6ꔯ~��wֳ]��A�4n��A]�������/��:���կ�@�^�~�)S�V�����L/���|���뇋���j0���|��_�:�(�@�_`{�3�I�y(+�k*�ZP�>�>X��<�b�'���|+l�nz�ƶ�q� ,UdC1������	ߜ�w66�\�x�/9!�Y�)�׍��̛*ᛄ��9�>��v��9 70��%��#����	xr,�YP䙔_��U� �k�d]RU,C�γ?�=��$�hK������?y&�L!K� \fcU���x}b�!R�m~f:B���F���z�o�_��G�%�F@��Td�C\�[$s�`���עy���6n1A�'���}���^�蹅��)��=�Y�C�f�����P�i1S�w���,�$�F���� ��L%�����
&G�3��=��N���D��.�S���O6OR�yx�x��󘸒��$w���9^ƿ�q<�&�i��KR��.n]��yq#�m�O=�����]}h0�veW,H<{��\C�sr����7�יV}��b��HYy9,�0)���,'ehG�X���Yh���520`!�9u�@���]98��-������O?�6
�(CL5����M�֋Pa��J��}'l�;DwY����yߟ}�zNډ����ɖ�׳�[گ�5z|�9y��/1t���딚� `�_+y��)2�om1�RF$}���U�9��#lw��Y�DIc,��>������Ѣ��6H�[2b{;E��H��nA�'�{F�)o_fį�q�������$�T��!F=��N����ff���ώ��Џ�by .�A.��I5�cƃF��t���CX��]�'/�}c"�"{B���}�	i�������ɚ��؄�MXX[�����LH#ksu�oL���P�8ÁߧO1�6Ap�M�\9OP7��ce���v�/��nn��]�lO�=l������Ht�Y�u��Ɵ�\�<hмͭ )H����3�L����@����V7�Я��I~�����P�2z���l�������$X[����g�B$�ǟ��ZS�؏���L�X�7�n�y̫2U�L�>��\W�:�fSI`6?�i#�r��Sh�3KI��mH���ͤź��诧�f4�w:��ف�r����m�0������P����q�(O����y#Ȼ����y����?��8��:2؃�Jy�=ol�EV3#�SNThgA/3��?[\���T�TLKAp�B~��)�`�NtEd���Yߔ>��!�"��fWn�(����.���Ȋ�ѺԹ��GG�d���r-��~��k�㝔�C��u;�%1��K1���x��V"��^����G�'�v�828����iD��IB\��M/���޵G�.�,"��tn�X7�.�x�b�P��I�Ŏ�ed~�D�Vg�j��J�G��,�)8���kʲV7��4���m�},6��1��0%>R�!�����eꂕ��Z��#5�K������Ԧ
��j�n��'3��":��	�9����L� sZ��x2�]a�׃e��R�w�����[�i��=Vv����o�"����1u����7�L��KŒ1}�]��eO7gZ7�����]�W>C����-Ӯӭ��ھچ>�/��ˉ�)�mR�HFF!�Vb�~ա����g�9r,/F&���s���ĉ�m�W�W�D�ȡ���
s�R|7���U�����ӋȟT����'Cf�4~eM��=�ƞ��?����u�R��1ۜ��6��Qg-�5шC�Q�C���a��5����gc[s�O��`�R��Ӯ]	3ӬC8I�ф�\B��9��q�+ʜ17G z���QE�2D���_]yM��T�JXA�!�geXw긚�Ewj%��|��6eI����������̧���o�� B���|i�y��v��w��XӼJu�8��i|��8�k�bc�>���WC�O�qR�'sTg��l�Hc�Ձ;��q�ۯ]7�a�}'���S<����5�M����}s0����Jz3r���ԗ�\7���N��� ����l�R4���gfԔu��Jg�����IA V|�	�[W�;�$qĚTK+��Q�/Dy���nBZ{�����w��Z+Ԇ�z��exS��m�J5,�{�zYB��5��1��eå��H����\F�K����a�K��O�ニL�<�O���{���ܼ�W>�3��E�_)��en���zW�GT�����t$=��>}*���6�S{Z+?Kp#�bw����xͷVL|�
jM�3T[�,�[%���|�k`��URjyF���ɫ��������n��@����P榺	�9VV�ܴ���c��xFB��+#�=4G^�\�~g�-�gv�A�����Q�&������WS&��'�-��'�l4=�AK���uok��ǫkc�ܚ3(]�zN)�u�����R>��}V����s�����&�0b_Io�����U�,28��J���[��1e����Ϫ��?�a�U�8��UEn@b�W��~c90�`$R��%�5��Ss�v�1�`���z������6��)j��6@���05:U��ij��Px/��{C"��ԛ@V�ƄJ�r�J�~��[)�jA'�k�b��Y���i����Ȼ�Қ�yZ>�܊L��٘�5��J�Y3�zi]J��!eED���M����
��k��X
W�6�
a+:f���߼d]J� l���؇��[�z��ՙ�5�?��3���?���[�^��l�m_"}�a�9Ⲍ�h3f��Z޵V��]���.@O_�����o��E��Ka������P��*���Z-�6��`ˬ���m!הI1-���,Z��-x9��n:���`S{��Wa���=�wz�o�w�Z�	�D\�&�	9�%jǓxg����c��O����&s��K��m�`�#I�,�/��=J�M���%�
�!��n�mu�:%z���E�{SJ��]�m<k$���Lz�����ٔ!��9��\r��.5��%��d�HBL��^�r׋��a���<5<�D��n�pv��������%p�$� �G��~.�N��~.�@e�g�8W��k��ɚ\t��?�)I���d���6��Z��]��4Abϯ����C_^�xw���+z��Hg0_=c�̇���u��SC ��z�P�06n�I��� �\��鿸�,��)ÊZ~=��RCR@����+5*�[_M�8����$E:{�A���P)�R`�{�+4�� Π����+V�X=-�o�<k;Ģ4�^��Z�L#�
��2���1W*v;������-^�Gf_ono������Z��.��^�4,T-��T'���!����SKoS�L]��뒛�.!��������wJ���)�zT��B����/��{F���w�Z��Z{�dW�ͺ}#�A��0&a����b�2�Ѓ�q�gJ����q�	('>#�YX����Kq�8�~������g����V4g�w�t��=�Ԝs��g婵K�wѠ6?���>3p%���NC��W�9���j��Rɇ=z�
o9��P~����A���/=��kP'(f������p4��Z+�fP�N-�L苼��峒�0�8=��H�����ȦSR�56���7�g�3�9x�X���48a��e��$�%�{o��j!���%�6�I�G��_5�~� "\:�O�i��*/�̗�v�w�~b���	�!�򦌀�f��a�$
-*�&N�85��&�i��]��k�R��;��_P��s�g��3Q�ꦾ���Z*Ka��S�Pcq�;��g��wecv���⚅ˍ^�׸�q��6_IL��b���e�ҡ�?ե�Ⱦ�׉�LHw�ٌ������_���Mv���߭�3��y�>Uf�|S��s��J��������4{h$�T�r�_��Z��{�Mv�h�a{�	�'5Kj�Բ�-�6	)�����ׂ��}�2��`Q����k��(���7�aF�k���2�o��z��7>���I� ��gm^$5%O�7d5ߞ���XpF{��Tx F]ߔ���2���wޝ���.A���ŏ������A�Z����}�Ҩ������I�G9پύ*X�'����=Eʍ�2*s(+�1�F꒙[��T��	J�EIZ�%ww�{�b9�s�P"mJ.n>ߕ0�M�A�rU�mO�(�����/����n/��5$�l?���8�q�������'������ ip;��_u��#��2��lGX&�a�ww�9�m$��~s�x�w�k ��ƒ4ʯ	AY�kBd���P"�pULz�|ؓ��į�������Đ6s��#-~e���Vs��eB�t^�U�?W&9����|�9�n�L������k"�=�~әZ�P1f*b��t|-��fX;%����i�J��{7���[.(����@��,W�4�kb%��t�0[�#�CM�����^ݑy�V}VljYGR7������ҫ\��2�$�z��gLԴ�'nH�V*
I�ʅ]��-�U�9i����ы:�2��r6g,��H*��e��"�dф QZ�����oJ�ۓ��z�B�"�#��ӷ2�ʰ�t{BgeWbWf.�x�«��ɑ�:k����l�^�R��M/ƃ�bJ��\F	)?��� ,�M��E|�*��/'�Ԉxnnv0�mpgOVļ絗��-�����^��R9����:�lQ໔�}�`��*q�w|�qG��sj��fblt5U�@��Y�߈�%u`�"��CÔh�_�% +��u�#�#_}���N��~U�
�`g9��X����Wt��2��p�0����v��G����ڧ�X{3�Q���FK��F6�bx`��⢖�8>>ْ�W��4L�\hs��a���c�tw�{u½���^�,�c�ƭ��#�a���#�!m�==>UT"��MB���Ms8'[�p����}	ótC嶧�=o�|�yMi��ߎa:��oU}8�#fO��VLac�GQ��lե���-_l���J�S�X-.�"�^�Z��������N�Ў�R�9�Y%�q��*���H�=q�A��A��9�n��z��m�-�ۉ��k��(S��у"WA)P����:�@��������_W�2p��;�le�+�����C�6uv�O*[	�و���,�w5x�o��}(FY-T��Q����-H����rV�L�$���.�[�k���N��C��Ȥ�l�m�>��ΡP��p��à,7P_����V���������q� 2L,�� ,|½��@����\���aΐ�$��AČ�8|[ڕ�$h�?6hޗ�^,˜�v徤�BmKn�!��|�Y�>)������:�X��nj֗�{;jZ�wE��U���|g��9���S�i�����t���e�1Ce���D�֊���z��I��v�D�ɛR��䫊E�r������
od��Hc]��I�$�O�^���Lx�{�ea���y��B��C�oӚ�9���=t�������#Fw��t�\tK��� ���Q������P�h:χ�,����P�;��R�ڑ4�ݩ����4�	o�A&��r����e��o����F��X�� �T<ol�>��M ����EK�<�쓊QJ1%�1
��r�3�}��.s9�<#����D�Ø��� +W������$�%P��'��w�^���pCޘ� �w+ ����`�9�qг�Η=)�=���y\	n�`[D�}AÜwa�����a@����	�J�>��y5-��s�sfZ����2/u��.S<t�[��h����`�����d_��ծ��ڈ����BF�.%2�
eAdY`Đ��>�(}��3����b��R�5��;w7��k-��uL�mk��$?h��h5ebM�>��O�T|o�Ƙ��+S���\=���d��#�7\&*˼��;�2��޶��S�q���θ4Yґ>�]&�w��s�T��<��z�|hG��tX��u�<Ay���������Vl5��<G�l�F�:�C��^H�8��w�V�0��O�/A����pUϳ(P�0����痤��
��˰B�&D�W���W�w����Ӵ�I�ɳ�o4�W,�ۦ$K�ֹ,�F*�m�*�a
o�&߀�>�/��4��"m3��峰oТ����޼�4�8鉽P�Fa�T���U�,ь]��?u�m��M�L}��X!-�]_�ˬR�����G�%E��{t���ց�ۣɅ��n�``e��MSp�MM\B�x��'rsfX2q��E�,��8�
S�f�y8��Ɲ�q������sؔ�Q�eI<:'_��Cw*0��v�`�l�y8�p���UK��r���:G
|����')<�L��ei�Dy4�X�(��.��"�#���a39HK�	%KH�f���H&�{?�^
��U��1�#-ށ��]E���|sP�H�wd�q�����/����.��y�� 4������]$�B�h����gQj�z�������D�W�*%[�w���{'�t�G2L-I/x��*��I�R�J^�F������~'�݆Q����FN�EH�,�C�`y�D�����:?��2� ��r
`5z��8j�qL]��{�t����/� V`��y���[�>��{�V��)�,�v	׷�l�(�Z��Jm��4��˽��[�nke��9��tc�t9Of_�}8T�N]|6�<��Ĉ������g�$�2 
���9�\�ݮ3���\��-:21�OV���O_B92,H�#��]~��������'�T�k�a��5r��s	��dy��O�sª�U�h2Dؤ9?��
�I�M~/���
d����uOcܻ��7��>~�&K��$��sצTP+M�d�ӺCO@ +&�?CYڙ[9^u�Z
�_eܒ/X{;���^�y����AP@l��~=���̳�N^-��'�,j/g�  �����Q&�A��&0ŗ�0s��Ҍ��!�!UҺ�k!�]J(P4�� �W��$�k��D��^���q�@�G�W(�u֩��� X�y���Z�Tb���I��Fh!1m!|���v����LZe�z��� ͑RI��S?hm7���huml�@/�UaF�I�������3Y!�7kM��0 }Lw�3��3�
(Yr���Z��\�l��f!m���V� 3��^����L���kX��
Ӯ�Zt�V,|ߊ�P�,.jU��iU-���sò�΢u�����7�<<�ME����@�8��@� ]��f"���
�����ʰ�I~V�ՏL�Ab��ͭe��l̋����YXҊ�$�{�zpT|�|Bg��E�3���$L=�Q׼�I_ma�Ν�E��v-�+�L��/,G�-�8�rD(�1�t��>�9S���i����5�Mȋ��Z��S�\����>㗄\YC�Y;c���YI������'= �G}���o���k�<�2�D��x xl���v�}:�(��-_��X�bql���̄mTJ�LJx�}la#�Xh9�	y�]��$7^&	�s�2�դ��y\MVc�\X��lH��)v��`���j��(�..˩9�js�I�bA�5ҐS�����ʞ���z��D����0�oL���(~�z3H������@"��u:�z�� ���)��L&���Ǟ8I;��m� ��B@%'w��+ep�W�4���ׄʍ>~/̦t�����P����u�u��y.x��wh|e��m|ᱧ�#��bR%�Lmq_�_�.�MM	�v��-�h�m��{F3`lh[��G�з��TT�ǈg�b��F����)�[�C��{c<V}�~�APS��Z�e�9����E�Kӽe�Ո��<��11�*_g���B������D�7�ʏp ����sqM�&g�� wJ=�ܴP���uj=o���S�jGw�g�ϻ[�����g z:Ee�p)��M%�Os�6�#;�-���§=��>�Vc&�l�=?�ޮ�p���4�����Юák���R͎�s��[���n��m!t�d���(���(Щ{��At��恀q�A��� A_�c������?N�U3��ZIq[Gi������5rv9���m�H�"eũ�q��c���`F��K����.�h�п~Hy�ҫEbL�ܩGM��Č�Q7^�����_ (3/<�O�����<�A���UB��1���q��g�����C7mKPP�K�y^�AЪF߬�����j9��R,t<��?^'��נ���V��[%��0�1�5(r ^I������-��yd��E�ۭy�G@��4j�5
d��.Ä���<��iσ�n��Kc��YF�AO�$�Z�����Xs_t��MB)�l�oZ�{q��hu俼Uλ�4�f��W�͉��_e�J��V�l���y4bj6�����1�S;�. )_Ӝ�?�[-�c�()Q �������?����������juA�y��~������^b3�!*�@P�y�g5���_�zϴ��u�� }ﲿb�w�󠬣��*2k�c�[�f#���~�4x-6��A��{2p<�@�^��E�zG��Sv���!�:��Z�\�����C�a�l�.����Ѣ���Y�`#��uVl�L�}�?�V�����i�A^�hs�b@e(�6�`j�Re)ܶ{riݣ���	:�b�h�՟@^�rs>��}v�T��]]�▬}���h-ڣ�����b �  j�%ѩ�ԡ�� J?a���IT<d��ۓZg>�gW�}��4.���/�:8���i�2�������������sc�^2������g��v�vt�����
u�mǌJ�۴<%z�p��vP�|U�/�t�p�HLm��~�Y�f9�;���k\;#T`�R�s��彘Բ&����Z��Hd`�KZ�`<����~s �hbg�4����86K�$,��&pK⣟ �-��_%D�Ѳ�*t�hj֫\���I�}#��p��pN�ը���^u�V0ף��S��u�7峒,��7r���3�-�֦v#�v�?\	�^�v<I��~*B���)�/K_��L���s=�sB�;��k���y��".���_��l�`�F$J/r��M��2�����TU�u��o۴�ɲ�ImV���ފ.'�(K��a]��d�|����:��X:��,��T��T�"��[�kd�ȍ���O������|�xm��o���`�i��'���O�4�^c���C�~�2띨�����?9�U��z,�s�Z#�9�
n�-h*�������q��,�@�8���Ԟ� �$n�A�(N�����/�r|"8ySp	U&�?�:&8;@]@CW1�ml��
"�xhxCLv����W6�n^&�䱣�*�]�����r������+��"��8���${��Sǌ����4��R�E�� z��[G�p��J��5���Ǹ�������IM���u�ƍ�_��4�i�{�v���]5����{��ߎo�.d���J`��X�]�;T�n���Ӱ�Lg����`D1Xh��Fׇ������CV���X[#��a�c0�}�kz���0o�sP(n�G��,��;�v��l�kDې��gʌ�Z���/2��Xn��ב�;��F�k}
_� �j��{`��Lo���x-�|r�_�VvL�[l�2�5qˠ^�F�z>4T\Y:�+�1P�0�t�Ռ�}�s�����W���qG�_�s�o|��ԥdv�V�z��Ӧ6�L�����q�+Z/�6L�Tڟ~�l��Q��!��\>�f�,���fi������>�S�p!VF���Ct�+���&�pj�,��+N���4�?��X��*Vg�>���3�->�t��	��m����Ҳ[q�G��S7�
Z�f�VQ���N-�+A��Ls$��k���[��Я���T�~u�Mo�:�i��!��Ib�ӧ]�=HC~VF]"[�� 0B�z��KM��M^�]I��ey����FuֈvU߬W��i.��)��8�_<����itpgoYD0����|Àv�;����Fb�d��a&(��1l�Z�tSJ�䷛���B��O����1��}{܊bX:m�T�q��^*
��Z�<$T�� �=3*�;�UwO��f�U.G:gy��z=\��c��qB�p��|�]�0mwڅW���T$J����&A���WY~���	���V�/G�}�7(Q�^_Uap����)��TtKݼ��	߭A3���Y���IH!��+��}9�
=��;үH�y��b��/ɨ2��\{�gQ$/��]�-�����<����������&MG8��L�GO���e�[��Q2Q�L�
p[���*1L�0�(��?5nS�ןH�@�ڎ�L�6�3�҉�{l�wk��`P�_T����]�g�B^
�>�\�W)�4���wz��X�g1��'�#O�n�� m5���n�������t����^T-gӵ˞�'���=�9m;�����%w:e����3� լ��3����f������Oq�S��ơ�Zf��I��k7���%�������F���T����u���3���6���;�@�e�)I��Ž�����X!cImpz�#���_��}���ş�+}n"!L���Y��a"�F(G ���-A���~����1,�O%��%P0/���� �A�[��n��SS�2{U�H�;*��l�!:,1	)�c�y'U��>w3�7�+e#L?n6�S3���ۧ��)���z+m+�	�b��)ݢ��1+\�v�.��b%�j��3�׿H�L��G��F�&u�Jiz}�A�dR[sYYK&�0�?����O��:���^�ב�p^yk���`���t�n��h
� �8�_Y ^	_?|�<�h(�w>��/{�}RЁXܴ}��#���2�q�J���*�M�P:�D�g�����E�m���za �n��uo!v��b�MA=N����c%Nm�TM<q 6O��؃�8Z"`��������Xw_X�R�[�S��Y�s>%~�(_�"�u�����)f�D�Ѯ:`��oPFϟ�q�AJzu�~��StXK<%C���kl-V�̇5�i���Y���V=�F��׿7*���tc-����j;\�0+rQ�Vo����m�������Be��K��fΑ5z��(�u�?��Ԕ��e���UD������+�_1��Ge���Q�D���ΰ���|��u��&�5ح��Q�T�2��bԚ��n!��/&^�o[�pU�_/�5`n9|�\E���⩵�?u�*�̃���0~�L�t�;�k�u�L�YJ�q�+B|�݈��	lw�����k97Sc�G��S�B/5�ba��p
z6���-ʦ���}I�X����GD
��~�F=�����9ь����*a5�ʄ�;J^Mז		k�C�p󌿯����ZMG�m��{��U ���feq9+���Ƹ��|��Sq�mI�V��Ζ�N^��Iܛ�!�(u��԰z)�ǫ����5�n-0�A��*Ә��k4ƻ>
tʆ���6>���\)�1`��	�%.}�+��̽(��ϸV&Iݩ�g�����&�KJ�ڻ��4/ �5��	-�`����&�/�'�γ�W�p42�?��.1�оp/ֶ{ٸzP(��qBn}1&K[ן��滞Y�Z��*�&���!f�/�H���h���#�$X�&@�����=b�7��P����/q.&�0�AKGH�GT۟Kd2�r�d*��,��Tf�fk��:�Kq�Pzظ���]�M�05�`���f]I���Γ,�X����AS���8�L�%�{���uw�>7%�2`gy[��k���ᱺ1^|��B�=�@J�-Q�~�ѣ�>S�ƴ�����V���p�,a��o�.��#$��l����N�բF%�*XNnk�n���Z/�[�S�)	���GS*��"��_�N�N�X�U]������1�YjBON7KBL����
,�Pwm�V�(B\���WL�o*�����~v�ʡ�(s*�C29Za�'@� u}���Je�h�W�<AQ��VZC��= !����vy<�֜9k��m]��iO��d��:څK ����}��/КP�X��6MГ�f+��՗ä��Bʳ^�+���)k�0;�׼�p�i�.����S:���h?�j��	Wܽ��j�R�������	Z�yiv�`t�PΕ):PrC��f�jw��t����G������R�BR������r�s8�=�NN*<�j�{sA���~�	Dtl^�DB�z �j��#�\<ܨ��,/jj#�$.;�h��G$M~�EL�(7yBul������aݤ��!�f�R��
��˷�3	��T/�����1���|ׯ@�}��Q.crx�����Nǃq�!!��lh��p��$iEDq�T����\�~���_�q�v���W"R~����_!S
1��D�(�Sn�{H�ӟ�܆���)蚲x��*0�kg�B���j�%���5�`>;#(�� ��E�[GE��}ã�(�GPA��.��T�K�CTPRIi�f�n�k���f(��70�9��}�k�,\�g��������{�"�����	HI;8A��yfa=Щ�Y$ku�6ZN���f:�T�,��^=9׍�ekїM�qBٿj}&�LV��ք�oi�4��{�>t�^i3qo�������E�Z�ߖ�v�ݠe�~�A&~�K�Ӂ"�@�_���g�r.�êY��a������h!%<������J�@��2���ӷ���B��d���T�܁F�8�he/
F@�ad��e�����Ѳ���Y�RtC��B@R8w4RZ&��)�`�l���޲�=���?�[�a���9&����j���K�����5�
�._�K��/����G9:Nbǩd�W��㬯p� �����JC*�v�0�9Csq����-��~@�Q`�C`�"�ʲ��%�K��,�6�=�v*�V"��"�i%�{�"�ŁP
�fA}�S��QhlL��}pLv��xӴ�zݎÅV��,�oQ��k��~;\o�
����o��
�P��K�����l��
�Q:�<n5�&�B���������<|ĕ�4�C?n ˅�i�
���������l_L�"G}5�4�ԠJs�����Ƿ_�3����a��	Q8��J_*��Mp��er|OR�z2���OS�+�6��Y B����:���ҽ*���cX³��*K�qՓ +���>}��]�PI���]c|<����%i ��sCI�r양�rG˘F()+�L�U�f��a�����T�ڊ��k�� ��O(�A��[���e/��o3����s�X�*�^�~��Z���u�d��x����^�����9*K�+��l�k�������wO�5��OV��eZ��D(���8>���?����kۣ~�%c �g2zw{��U0�-��2띴�کP%�h)�.�2[����ݠ��rn��c{��n�5�2�mɤԧN�d�,�z����W !2`�w,�Z�z�],���s���]�T�hu�p{�h��LpI#�y��`�::�B2�5��<w�	��'dg��y���f�>&�:M��+��M�g�Jz����y�+U�X|��|�f7�{cY&�Co0嫥��2Ն���7m��r�L������@���+���`����*2=Y�R�s/��[�\����]y���2�$����%r�\�8�C��{]4�����_��.����Tl��E�?�t��kRT����M9��QT�٠��ց�9l`d}S���3�&)uF~;��f�s棓�8�~�j]ʝ�,r)L������ƞ6���5���ƮR�˫sG��W��P,]m� ��$W̿#B��"���H|�4�l|B��'��>��f7�G�+�S��d�z�+l+v�V��Zb`�i3Υ_����]���_��ת0[���:]��3�~�X�1K�7Ɩ�j���'�e�(��/3�Y��q��J�-Ixٝ�,*�Ƨ�`�$���c+��#�Z'@k�,!�az[,}`KT�E�nXQ����x�-&Ma�Y%���̓Zs�4v���,��̍(rV�5N%gؓY�5M��!ߜڛs��{�q�-ľ|���D%Ax�O�<׿�������w]5qK���q4�eTdW��gʆv�hޱ�����&��$y+m=B�yػ��h�qiFR}Z��xA����5�_� ��9��Y��g}{N���̢��ʊ��i��X�i��pt5rl�In�?x(/@u���:|����!�}�W�[y�Lbg�/Wxk%�w�����̚�,a����-S��.0��tR�]�;��S�\�D�"J�ܩ�Mv��؍�����I$.
���rdؖ�q��$�{�25�b��KG,���r��q+��3��<�fX��^1�L��|�O.�
�mq���J�6�2ލO�SA>E-,��F�-�~|�q����.)P)[ٳz����D!@f����m]���  ��i'`D:z���k�D}��a���prF�h��<����/��|��'�I�+N�DSؽ���Ʒ+�Li���!����۽)<���^'�
%��ɝ�yǎ3��O�P������P�'�Jn�Š���&YvjQ�c+}���T�sp	��:�������6����-yr���8/B����-�0PG){ �C�5fɛl!���+��vګ�j&"��|�����#��K���#Z�y���i�L�W��� ��t�5\�y�i�K����n �j7���� �ѧ�ӧ���ܘ���d�'�x�f��$�P�{S�"�X�#5A"h>@���z�����T��(���R�vv�L)�lٽ�d�$�.k�3.!���(��.`�c���X:{l)%������ӎz2���޲T4�#U#i#"��?:*=,��aj ���G*6��:��51G<S�
Ƴ�7�WI�^vJO���+ը\���9	8JwĿ)���p{������,p�	c��v��j*�,ٷs�M�=�y�5�M=�.��.n�6��ql��-�Oo4Y� \Ĺu�,7[~<z?J�&�� ��
Nh�AJ��\v�̦Z<�;�8���]Ł��@�[ۻ�
����ӓ�i�\���1�ffi䡻��`�(7�,�OD��l��썹� �v&k���L��g�h>�3z�����U�#K���;�B�W	�5�&��Q�1��S54��,�3<Ogx>��!�6�m�?�=�L$��鶔5>{�Ǝv��(/f;�b�Ł�+�xA�q�/Td}*�ZH|�<X�	?�a>�z��N�c��~q��%O����&C�0^Q�N8�	
td!������PH5N&���q&��ᏪFU	�&�XS�jZj�H�ko����.}&I*���!MjQح	y�:��&�a`�l�,�1��G���d���4S1,,TJ��	�*E!����&�J�"�E�NF����P�S��%	5��7�v�Ŋ"ڢg����6�ǡ�y��˒_Y�t-����6ˣ˨�(>�pE��G�7Cw�-�����[b�*ܧG���3����;>%�MA�(z�I��/�E��P��|qP�}=�I�9��ҥx�!�X�[U�On��ѭz�gK{j�P��U��Ðwg}�qɝ>:�Ď�8{}Nx��N
��� F8�8�ꚨ��(=�Q��u�$� ���+���~YG�����#���ߵ�w8`�4��5SҒ���c��׾���u�"MJ�0����!�.�nȇ� �Y�^1�/�G��y��^��8���w#��ӹ��T�;��ϙ���dE﯌���ȅs
XTНB�u�l���/dq�zi����فI@��͛O-)�Px�W�P�4��[�K-��i�?7��_�TUBp\��N ����$��(>)]��m�0]%�,;���SE�R�Y$�G����T8u�'��f��(�fĐ��mGL�5�01��}Z��f/jxw^zȼ�$@�|x!:>�č!�f�O�z*�L���3�q��N�!sy �*z�	{�Y#͡:�u����<�,k�+�>kmԭ��7��2/�#������.�s#ObA�6��o@�.,�E{��1[ �f�YXO��ɖ֨��Aw��Ŭ�#<p���W�R�s����A�9�قKL,��NE .!�l��w@x抭����Ԟ�(>r��s �爙�� ��8q����\9j#�{6͚���2�z XZ�斛���_�L��M x(���xo��@������W6�Tp�6K�Iܢ۟��Z�BJi0Ӆ�ղ��"tֺ:��<�ϓ81�?������"3�ݚ��uKCeMI��*����N������>YZ�2V�?����N�%� <����VO��)��N	�7��S���p3�����q�L<s���G��r����^���`Y����|��i��yX|��C���(P���O�|�\�Ê:6��ѭ$v���e��6H(�d2~�u�Bz[,��QU� �B
��*$�a���n?̷=�0�%; �f��74�E��d8@�Lm��}�N?��k.xRT�HsX:��1/^�XR.�mz�.C����;"G?�E�Nx�C��Y@b-�%�p��oŐ����a3T�J��� `�!^(�\����½��Ul�����mȱB��q6�n���P��X:�	���B�U;�/F� ;f�*�c��}޺��𱒜�5d���8���8����&;)�CY/���q ���
~oki#��8�X_����M��F5z�j��3y��g���{��]QU5���kM��d�Z���m��?B; �@���={�8|�"G3B	&�\�_�q9	�ڧ룸'�X�^J_�����U>��7+8E9�Zk�/��>b6H�m�]��=G�M���O�z��JӔ/��=��7��`�}13�ؖ�*<���0h._֜�"D4��H�O�병<�-+ ��[�s��Q�N ,L~j�2[�"��58�M4G�׈���Bl��>%���ӭc�^�_J'rd��ۭ����6jQ��H6���G��,J����`���fg��F<��ī��Z�R���&�+�\���&�9�
j����<,I��s�o��N������ڭ�(|����޽
�������~���Q�Y<_��պPb��h ���ص Gzh�Tqf�\�)��\��a!�n����G:�h��守iD��������Z(��(��*z/����:�?u"5�:���$'ݓM�p��k��UN�w��>e�H̀��r2,���0���P�vl�]C�}��vyB�iz����`/or&�7[�y:hwS�y�Ez!*�\N�dU�ܗ�o^&��,��~5G�ァ�ݽ���Bi��i�Ç���M�ʞ��|�Օ�����JS���}R,�Te,v*^�R�D�a��^V/������֥I����+s!:*ʳ�-\�3@I�6Ә��ЍzvwO��>]z"�y���{��z��h��:w�na�S橣��x��Jck��D�S�x���d�����+}U�Sq(��3����R�6�q)liE/����p�VZcܺU�OaǑX?�Z���k� j�2�08U&0���j�O �p�*��}p��̣Q����Fk���W-2O@�H<3}����Zޖ��{��O�),V^���wy�j���Îp f8MPVv%K(�E�2�tI�`��c��I�����p�Hdn�#�ي����4k@kN��z28'����Ie£��� ���Zah��I ������=�}�i�.�� δZq��T�E�i���iO�L�t.�h�H��eqz)C�l�.��t`n:L��X*�TE֙aH�8��M�*ѡmi��ӕŅ̷��jd��@����\��D�%S�4�ſ�z�����CR�����$�O�.<}�q�Q���8�K��<��}[��QC���d��\�80Z=�F]��G/#;�׾�ح�8�30.0������v�'��3�2n�t��V����+�p��.'P�Acf��DPrr�+2�D��'��z�!����S��.vKRBpyHn���:U���-D�A���wu�h�i�n]V�|���z���A1���WZs�������o6��ѐg�"|���.��jY����B�A�y�~��N���ϱ�CEs��~"�@y��?��L%��\��T��*��w,�f�D��)J
����� �<��
S.�M��85�:-�ХD�7�9��R��W�� �w����L��p��I�}�
+Vחɫ�g�b��נ!2ܒ~uw�bv[�bG���qN����s~i�W��jD���G���_��ò@�b�~F��}����r�ۧ=�#:�%"׍�g��L'�����c��b�u��x�7�_�
�47�PIZ~�]�`�*��R�co��P�*b�wO4����a���#�)Mv���;�k{�fzU�k˜�ᬭ���!�|�S��������f�v��c���h(C��������j���Җ�����퇿n� �C�-Ȼ�_�k�hsŷ�b��#�U)��-Aq0� ɽA�#J}�1r���=���@�u��)2F|����h}'�/{��)�_������Hb�a� ���X���� �]���d��r���I.S��1`>��r���*��^�Px�ƚT����| )3;�/��O�N��+����*홑C%L�h�|�z���ik��<�W����r�Z^�=氁|H���R��a���?���~G��C$�_ߥ�Q����\�9s�%ǅ�Z3�~S0eUG��۹//`�[�������E�ݯ��|��S�#|v���iKS '$Ee�A��h�K�#�-��!.�C��¯�t���E�,?���=�W4��>��R
����RI�b����R�epB���K��)�����Z�w ���
S�-��l��N�,�
ue�難��20~���a�e�`���$�^"L���T���������a @��

�ឩ�w�hd���M������!/���s�?^S��P08��\[��r���Z�}߼M��|
����q���RdnY"�[q@��q��T�������B�Ru9��x���J��y��v ��/v���ԖP�\�B��� �t���Tyj�b~Lw~ORm��2�z<ų��e$��� � iW��c��I�V6��A���Y�R�4��%,�A�Χ��6�Zs�~���K,y�}�]+�a��Y�& �̷Z?4�W����$h�x���N��!wG�c�Ɓ�H{C}eT%�}��R���n�I�[,α�9�<��K0�@Si@\||WC�i�s��d���j��Sa��E,	�ʼ��v�'���Y��}yq�>�M!d+y#P@7��s��T���%���X<V3"��z����4�A�P<��q-����o�6)����>�|��|�ф<������їp���b�	��-a4�SX)�}-晢�(t���m��Ed�P4�	9f���eK(|RL����bĔ���F�]W�ࢧ;�}#�-a���	ҊoŘOwNލsh�?4j:V̟Pb��`��P�y�+c�b���H[��'��}�\���NKi�4)��F~�$����z�̟'Š��c���l�{�����:=�p���N;q���,5��0��p�OL� �L�y��������!%v3����kSV�g�I{��ʰ	���u-N�3���j,��O�M�,����9�$�X2q��+���h���9�Z���l�ՠ�{W�Cb�\?Lw���nd��!_����ً�ڻ�d�.���G���X��Cf���aӝ���k����S=W�y2<��7�J����vcG=z�������Ԛ�Q1���%`����c+}{~7�6=��Ge��+��_��o�(�r�rS̰!�y�6�����b�,c�p���|��«�ˀ;xh�щ���Y�6Ou�E�-�ͽ��(�� �����:X�4��%���i_�|r$���7�Q����D�T��6jnK�*S�Z��;݊��= �y�֯�X�+w�ͻ �#��={p/cz5�oXiN��@����_��d�D~=*�=�%����ɩ	.9$HK��}��/֤�l\�5`lǪ��Q�9jڏ�f+CrP~3�o�]bsQ��y\�gQ�ف6�5��I#Ji��cY�VC�ʱ�Z��Z�lFӜ� \kuc�\�����wT�n]�׼�z�W2�T=���ϵ=e�؈�F�-�`�S�[�L�.w8g4:���<����O���ܴ�0,�Q��D'�fB)�e0_��*EEEB����9�YSmg��c@���xQ������y��*�D�����P��&$_����L���L!�J\<�B,/����]1W�Co����2���nT��C!'ޜE��b��-��b�U)�%�.ӌ���)1�h�FR�~M�y��(�b9-S^�v��O�A��_v�T	������{�2�l#5�����B���˓=�^�丌���Z@��S_˥�eg�o���_}�-p����|$�>����<I�K�7���k�he��&_��{�!А�Y�xa�iU��2 wC��;b>�r�s����Le��-��ݓ�y�(�_�e�� e�L-�TnH�����z�ד���
aE�,��k��n""�FA
̓p-���?1�_��(�9�r1w��i� W�Q�`Z�Į]s� ��E���\� *)�B5 ���C�h.�$����l�\�4O������E�EI�Eb���8͹'=�'HE����"Z&3�&�ёbS !@n/�@���t�
J,~���f- ����u�� �z��f@ڗ�nsqg�c�2��� s�������+��TtM]CE��������a�λkFS;j\R�+�HIW���>�%Y�b!�m������z�M,�c�^��N3��B(h���ʹQ�Y���~s/S�&�S�=Uh[�I;z� we�g�ف{>�ҲO(.��T�*u{����ϙ�yj�Y��2`�B�>�&�R�ck׶��sX�TliA E�P���S}Z(
8��4砄����<-�c_�|<Y��%����G��T]��؅uǡgpd��ݧU�E�wjc��'�ι����#a�<��X�'�$XN�&�4�8�[� �X���n#������rEm�_[I���3�t"KU@�6R��]������n�HI�8�0`�|�q6~.��[�8�O���VF�c�ae�RT2�jh�7���\�0��uf̀���e�u7�ϗ��A�t���ւ�+�pR$�ʥĐ^��A��9��t���\�{�2�h�G�Luv��2�/^ty=߲l�'!X:������׊���H�U%oW.�n�=Г<X��nUQ(��*^tٴ��J�༼��Fe��W�08ja�y��O�K.-�;����s�N�� ��Ԯm�?Z��}�2���A���<u_�su�0XxH/@P�nZn��ӥ<t��{>Hr|W�@�0��nH�nxOo���>����(�����TwiƗl\��O2���֕m�B���gX�:w��l��D�|��D�zd�I�4�V���&���H��O�$�yZ^<Bo(���g�����\��@ة�=����p�J��O�T��2ܪ��V����N���E�RY �/�ٿ ;;�fou�^�z���bkK��N25;;�	�X3�U���#�5�+`ܱ5��+�W���F
�7��Q�Zۘ���7ߕ�Yb��N>Nt;�\�r�u��HL�zU\��,�<f�@0��=Y�δ�r�I��|,���)��L �8�9� ��⤰�����1�Fw�"��I���5ϔ�P�-��K6�T�u��X79���&��U��U3�O�VcPn�ٟ�۟�@��w�VQ�;���sz�XX�R�-�F�5;ީ��t�_��C���nF��/��|ѕ�=ةe�^�w�D������?O Ǳ�/W���%��!�ð��~ �o8����:[c.=�}KG����h<̈���t^Fq�c�����"w�c�[KY��/����������s�'�iD=����Sy�Q^9�n2M��сJ���������m����>S�.QZsY	����,G��֊�|�;b�=]-���T�b[�0��0�RX�ʰ�A��ی��޾w����\%ɲ�')���7�
��@�&-/����6O���Kv H�xR��o�\S�1ބJk��}��B^�L��Y�Th�騰�'�'�dMi���Wʐ(u��&�$���JS�fJ�ҝG�����SYLe� �T[��s0t��C4a��vw_�m��!˂��W �`Gi%7�2dQl����ԉ$����@���Cko�z�șy�s����W�b��~��;n��3��� �ߥ����L��ô���X�!�I%�3�8{�1]M��.�|C��O�@~e�B��I0����ed`��Ȟ)�b���88����QӼ��~�QN��n5�ޝ�ThA�(RV�,��^�qP���W���R'?58LS V��"��@���Hgb�O'M��RȠ��+�yY����:k�Ļ�~js����Ȧ�su�;�v�ف�l�3<�}�yi���*�:�*b�i�d���p:�ȷ�'��$���U;�|����T64LC@�g�8{5�=_��h�E/�JB�u�������=����G>V�j"}Z�.xG`oD�-m+
t$#���������S�>��>y1����dLR��|>���<�#T���h�H �	�����~�ӧ蕈�2��%�j��/3Ŝ����0�yŪ٪�c��4'1۷�n�61*�,��i��c8�A"�v��p�����2���EW�
���G��bB��C�;�����	: ��Ju�����x���G��FA"��i�z��wN��zNN�g�fo��
���-|U����6�g��Xr�⃮qCc����~r]��i��<p���<� Ή��:��S��nټ�o�6 ArE�� ��I�M�?Dh>�T\f�S���)9!Y\D#ra��dy����|o�#�R�:�Rj�3q�E�	ъ(�gY�BIW��!!\y�	�PV�6���6���MZ���Y�R�J7$eb�Kx�4�q)b0tK�bc�d6]9�{n�g�ơRG���W�t��/���IL4����I�3�lf����W@��ϴ9�GWkx<�I�����:k`��0��О�{�2���m�W������P��� 5��>Ԙ�;��SMa�u���O���0��޴�}xݶ�� ˺u����[��L��q����$�|���71bc�Ů��x��x�#���n��O�8֛`�?y����^Z�����L�$u������q������7|_����\�Ƣ��(�I����+�~��R�6#k.�s���qC����>�F�ܬ�g�F�G{�;?�,�v"�	9hdÖ+@O@l�U!�R�\�>�7���c��J�}[Ǜ��{����;�Иj�P���[̲��I�.�!  hLԒM�r�)�Ch�O��PȋN\H�i���l�T�qF�8��+~����L+c�����/+|z�
D@�U�P"�`�=~X�4�(�)���r5�}� j�:��*=��U����QI�>���G�~��
��b�Ο�)`o�ħ�[�μ_����p�LC�36��N�h��58�(�x�ڕ5�peq�ݪ5v}�4 0��^=0)�F])5���絿��db��������+��u��Qx��Vf)~W��4#U0F��te�p�J:�6��f�K�Tf�H�;�\�����b-�b�6�K�#� ��nF,���٪�p�m{[�e ��q��s-�M�^#�Q����g��ϧj�n�U?>5��Rl��	�4FO�ᵵʪ��M���KŢ�L��^�2]�T'ya��9�,`}'��8���E�3w<���T���W�V8��rXG� ��/Іve�Sz*��5�N�x���q��(�N�*{��Ry��M�%	�{�E����P�78�����G.C�r�g��(�{�	TH��
`���]����{̕U���5D
��DRr"�+Dz����w"��?��5�G��Gk�Q���u}���^��}UX�����q���R;�iI��9�xhB�D�&4��'G�EG�*�'��N��L��'�+���;BdR�D**Gu8���EHN��]���?��}|3��x��Q���I$f8�V�	���	�}���x9��a�����q�Mh�E���"�f�钔*��Y����
݅=ۢ_S���):wL�֪���ejD�~�d{��~t��������l�)p���li��Z՛����-�T�3�_�	d'`��R�˞J3����I)|�-�c�I����������/R�q�s�����B����N�Y*�N��_O�b�������?�I�~�1RY��� ����m`��g,4g��}�0t�謙}R���n��]sYb��n�,���CD�H�r0_������ɛO��]��B��u3���k�s��s���3����Ƚ����P	����Z$�T�Nі���T-����C�L�#Ϭh�G:L2�$�b@=CJ�}�v���V��˜��Ψ��,G��?��pv	h�����߷s)l8�z̢��P��y|��~74�-�k�e|G;[���W�x��z��KGC?fQ�"r2�
�R�n�-�R�m���f �����= T�|=R��%黅Gԉ�b�֊H,�1���ق4�������sJ�",7�uDh���j;áZ<�B�@�3�W�#M�h{P�E+� �V�l�N$1���,ӰNq�m��A��x0��;WY5��{��ʨ"����Ș�L�DP���U�s���J�(+�PV�=�C�b���˯<yX-��-ĘuKz��te.�((�&>���{)��K{1Io{#�0,S޲h��� d�o'�� ���$�ƀm`�����!�'F��;I� +Ņ��~nS�bZ�5��(�ڟ�.j�Q����?g�	V�ϫ�[p����"�3��_����"���v�J0�]��Q�w�t���9	�W%v��#�(�/Ei&�q��)�i����0Dȧ������aO�3�8���۲M���[�r�;�������L��<�|�4ϧ�Y�}I�jօ���Z���Ή�� ɽ��+��UI=mͻ�o�^���������l�r�g������\�ԅ�ۜ�L�S�0Y�SIl;� ��O=�p�T�vǞT���rph��OAf^B��4l�Ot�t�?L�M�Wa�2�"�Z+`�a��}���4����v:8�cA3�����V_��gfg��2�:���"�m��qꙎ/U�� �6g�I�ڏ��锇ʿ���$�j�T�vntt�v�3��:D�5��-�XI��\I���C��E��N��B2���%�]!�J1�rN�슥mb�%�~I���0�Y?Q4mm�Z�]�^�fbz�d��F�ٷN*��.�N����]i�h:74\џ��}���g�6�Pa����;��1;/��LR30���x
�?�T�E k� h),z4L��Zǵ���=/?^k�I��>�;٢Ƞ(�f`h��
�A�u�2K̆�K�DEEÞP��P�3\'h]�� ?l��>�μK4��[�z<�o���V��X=�|q��z�h���������g��xR��q����n�_-���E��q}��4�2#�Z�#��eK{=�h��=@|Ɇ�Q�S|�P��|�\T�u�����i-�vp(�n�	�gRcȭzfw�{؟+�-^�E��kʹ�||���8ǉsv�e���|��{��9Q�f�� ��I}���%��Uʃ|�s-���l1�p���w_�d䶱��8���F`�K�AO�u�ΰ�?y#��ܜ�`���,ex��h���hkn�� 距�JdK~�2��t_����|Y�
l��|��v��!!���������?�3<l�?�!a6D4��&x'DF0���Y$�wp0=-�9S2C�������ɫWihlD��̭M�����x�.W�԰�<,Gon҇4�����cn>�JN�#�ȶ��O^�I��W����
"V�'r�'�"�,y?@e?	)����XU�D%YŸ�Qp�ؓܐ6�H��qJ�_��l��[1t�:�ͼ�+;�lt�v�v\! ��M����!�F	cǽ��2t���`���8�����Y��r#�/w�Ō���q��Ź,Gڇ���j��	�F�/��V����;�/�ˀ�|�Ds {O���-@��h㮖��k�xR��R3�r~��W�.I�4���{��i�'�=�iX�`Z���=��LUT�Hc.�:{A�.������ׄ�l���^�U�r����W�7�M��2�J��z/|YZ��F��h4h��
�\�2�GU��V�j�"RRRi,,,2<�Č���	lw���;� L�v�>鈑�H
����?�z4��h��֘�d ��b���L������&�m�3f>-)?�*��٠�W��ܜ����ν�Y`5G�K�z�xC2�-J�nE�OM�a��5adj�е�w��7�Ae����)���|�X-^/2�}�П}�QV�G�(B���q�b��6޿�f��{moC�����]���R�ߧ�!�V��R��_yfcl>��,S��}��g�x�D"-��8����l.����x�귆�B�\���.�<�}����/�&�T���t
pg����LLL����#�H�q[H���.z���gT�:�ҥ�1
��]kW �"~WRb��}�9_��3S�����.�Wy^�劖�����Y��y��ҥ���n$�U����J�6ЈQQQD�;+**��{�Z$�������
��#�����!g�)�ħo��%���$麂�Z:�hO�÷:^V��H"�Vu� Ӕ��5[�R�����@]��`5"`�!ӻ�X���n�8�4����?[����8��L5���V��n����������%f����t�#�AL(^7�C!pk�sQ��c�z������S'�"��^�FD��塎���W?�.��c�q�p��{�o�׮Sy���i�@x�*ig.��GOV�7�E^�Nƕ~�&�Q��)�p�q��������T��&777�"4|�J�'65X���j?ʻH{���Y�e�xWkM�n�����_�p� $����!�`0��,���}gº.0��kO�V	��̱�-tV��$�[/*�J4F��Y�ս-J0&��M�i�p\���+��Jy���! +�:����P�T:r9-�^�l0���ɖG������;���׶��*$W��H��qwX�E�1Ͽ��J��1��X�j��K�{�(-�ݹ��?���C��ф���gJ��� �UN��_���lsqh^
yJ#tC=5D.}��3BZiʽ9���������3�r��"��^Z"�F 
��.fH9�*A�-���މ�x,��g��Vjv <D��4�������*=�'��;蜼63u���EIFn�����W_����`oK椧AM��}���h�x��C��g��V-ti��.P�8[����B �'TUU�������X��>`ͧp��C��!��F[�$����?�R)Ӧ��6U*:��:�ӧ[9e�<Y������.�]����%�t�k���`bN����]B���O��E��/�Y�Z���L�S�\�~����r�lÐa|,8�Q���?��z�N�=�3F����Uɚ�yMS�&0��
0�(
��_�~��1��*:c��4�62&�4	eM�B�)��7��S�iqd
i�R�������:�yԹS�d}��sr���m�bP�'6zed�1]�I4_��vRTS#��q��%w`��|$/�_BQ�7����gHV�8��f`��Y�!���I �t�{*�'���iB���"�'M���g:K}q�l̷�ׁT : �G��e;˕��Y������!�вWR3^�_��|���=k�/-�z ��ے�����2g[|�{<���kk;�����&����&�z߼/X5�;ԩƆ�=����n���615�i-�/]�Ѝ�.M��jc�#��}w5��:�������'�T�_�&��v]4�:��L�;�`�̤�O��Zo�nL�� #��|�>95!�FN�Lԡ����6n�Wv2�u���1���C���y0���m�,�V&�P�����z����n\*L*.�\��>388�W���e��{{���T[� E�q�m!�R���ZqQ�a��,����j�~��e����7�s�7�w�@w&[|��r5$~��q Y�}�E���e���QaF�ncUNV٥4\A�Ɩ��u�0�-""bUO�����Jz�w�Η�6\���Б�N]���շ�u߿��erV�" �#%B�Lgw��0��r��W=����{%R\����^��O)$0.d�7�:��l�-RNA!�����I�ko{zz���4���f����#��(�J��� Tt�GƄ5F��}�	��Gcyi�?��Vio��Z���
��9Y�����4��yGi@�7&,�K=4�};=��ߵWm"M'����Qh9�D���c<���u�����1Wܑ�m2(<~��Qz���M5�$%$��i������oՂ�̵�K�i 	J�=j�����A�8�*4l$�����@�e�x�0~�1߉z��#"Ybb+׵�xP�����	�ZX��Ht�J*y�@$��z�t^
�mZ��xA  �!����J*Z)#c� �iX��^-��s��`�]D��������z�]�44��ñ��Cn��I�9��Վ���^ /����a�o��`�l�z��6)H�/?���f����z'-�o$�ɭ���R#��
1�rphz�����L����g��7�f~�% ��u����X��������I(�[��.�f\��wƶ�}}}n�;ȝ#�<-����Qy��РZl��J�ų=:�z�E��Lrb�Y�������Ttt(!��;g^x�ޟ����HyFV<C�K�b���%!Lw�D���s�Ѵ�r^P� �T�޽�!`�ehx�c�/���an��i��GNS�O���Ó=,o�dO	귄:�7!t�.��&D�֣j$���y���J��Ptp�l�yyw[Z[	#q���6��[���w��!X],��Ȏ/R<�,r�j:L�S2�V��m���<�������N�!�~��WPP �;444����Y�s�F�^���~������t��KJ��!jg���;GHS��V(��o\]���P��5���Wg��KKgdg�����̯C�	�%���*WF(�6���ޟU̒TS���q]t��Z�+,�/tFq2�H~|߂��q����5��񇌁��R8Q�cz�S����v5
���)��xy���:����1�0|͢�&�������fm1��a�!	ߥ�
@y�V;����^�ם��@���
��溍$��C8�4�K|]�BM\���o` |����Ռ�Q��EC?�yϛ�-;�F� SRR�@0EA����L�����2��p�Êi%?��n�!���!��}5%Bx��b�����ɷT�O��d��������z��F+8�І�Q�aaaY��؇��X�|�_1�c``�.��d�r��^��.P8�%��������Ei���|A
bLղOKs5�� �8Z�\�F�� �
��?d�Ks�7�,tl4���]�I��7�ފn�_� "`��w�̓�xGlO�Xh9�-D���6��uK�Է�k;쬤�4Z�l��k$' N��lqq�h�6��Ҭ����	M�!��65�����(�L[����㝩����֏D�xPa����:�\N;�05���GI�f��V�tyF��\�95�#�8���@�K��>�s��+�;�����)�I��d�rs�cKV����Z����a^.��m�r%�B+�a�j�sii�[�����W �6���.2���=���l��RaIq"��;�G�O��x~�58�d+"�%�U��? hM�M���볝A&������y���+r��o�O��f-˺��P���UD��Fo��k�=����p,3s��Wܨ���˳���W�lI��
��0-�U�p~�8i�Lg||�P}���恣��1pq���Z}s�$��[Z[g�wS���%��;+��s�w�-�;bڥ��R�N7�,}�Y�X�:v���8�����ӹs�׏�+�����,���箋h�1Z���Q��'im�y�t�uZ��C��qCI'��=<&������-��*i��4�gҰf�L#�����@B�����ўX$����R��ܷc�߾47�3{�I��u5{r��AߟS��ZiIC����TEho7����q����_��kw�i)��N�f�������k��W}��HQ��R��⥉tiB(�	=� �NP�R���AzQ ��[$�WCI��?'��_�b)�0sΞ]�g�=3.=�Qt�!dwx-����P��{r5��"��j�|�AX����Yj�������kV���k�e�),X_`�Z4Ғ��ѐ��t���ĝ�`�^�����ƾ	V�����_��2��j��>:
��Ž;1�6���V=�\�ճ�G+� �5a�e��Y]]]k�������c���1�7 E��0��*@�gK�e�"h���_�
G�4�4�
�����Wbz+����P���:ry�9�������7u_n�f�	�H�L"���v-������1(((�S3Lz�� ~�<�c��oXj�������r����yS�|�=f�*�����k���/�l��7�9�W��^(Wc�&�U��#�+�����`o7!��46�̵��w}�����pU���L������xP���*-���!��,�%���`U�C[�v�~�p�"��<��^s��3%���[PO8�^�{٩����/��<�ޟ^�k�Ř�z��S�f_�����]oy{\lz8�/:�:-]zQ�|}:55!T���ƖY�Gy�A�=�C��+�ڔ�i�Q��	�lO̮����M�m��>�lK�_�P�Y��+�J��5�܂���3N���GX�h�)o����<C#҅�X����b�go��˗!AɖC��ۛ5��嗩g��uI�}�x�����YO��a�L�7�4*�4�LA⿂�7�����,�`f_�PW�ќ�b�����2�OF�>��- Z_KI�d�>9�a�j���H}y��!$���+O�0���N��A�۲��0�p42A,WVnoM�+-��зρ¨-�q��9�d�����M9`��-�����
O��o/Pt�F^���m圣ߴLX�52�,��e�k���Z��:z.F�iatA�4�z �Sz*��?��r�]�)���@�Ԟ�~���ߣ�m��%�����ޮ����f�/; �#��e�������2�a���o�^{x,��΅<P�n��a{��~���&�\P7�������H������)8�*�LsJ�鱺S�~YsH���K�k�!1uw�i��n�ѵS��_𳷺NgU-9����AMAM e��U]ӥO�Ԓ���P[���V�����M��N3?ۉ���>}��*+ua���+y�ֶ���h����kc��nY�Fvn�f�-�Llf��+�7�����^� ��v�����_:�p���bO�!|"oG���t���{�M�C'�qg�-�p�m��kB.�}�u�����</�R�,s��0�o��T%�� /Z1���L��VJ�!�`u1W���U���`Y�b��]`�_.�a[��o����5# Ă��	�G�bw��.C�6��8L��MFM�y��&&� �TH-�h�ͽ*&��!��ÙL͢������Y�n��:�u}�ׄ��RZ�4�, "�u,T�55��ĆR������_Ň[�h����9Q�C�\�wP�w�c������:<����|�t������B�����[��� �N�_������c����K��=STYfi׭�X��jv:�z�r)M:���tz�!��lU�A�÷����.[�v���e��k���84�0lU�0��穝ƴ���?d�A��
�tH`�(�_����튒4�I��k�� :rb�ѷ�ǽY�H�L� ��e&����|d!��.
�p���J�ysWˮ��PY��Px���P/���Kq_n��~3@n��~N��pM6�#+g{�[ʝ�%kS�+^�t'�4F*�?4��1ʠ)�w�c����!:��� �yI�0LA� �x�K�Q\�.����Т��b%��������p�6y�`v_�R�ߦs����V�5;D�,'t��]! ��FV��D5���p�0�/4����fQ���+�@��M�A�
�[�x�iS��2ɾл�RQ��(zѱ}LD���D�Cs����� ϩ�mhg1����T���hy�׋�L`��_n�k�Y�0����S�k��e�����:K��?��4珔$�F5;0�/���2��PG2�L�ݓJ�����*?����dz����cA��ThX�R7�VD\\���锝��R�ؿ��N��7�Z4C��p��W���j����Y>`��;�{GEE�i�-��݋� ����6ճt��~�~��l�ĩ�[o���`57dr)X�5��2���� �!��J�܍����]�C�$�����iW�����q�^���zp��co�e�(������*q�R1g'M��+v�ۊ��3|����yNj�^���U�������M��\ܖ��i���޻��+!�?�b�ʰ�����
�e�T��0������P7U�PԀXT�����N�q�{�a��EipL������)��m�̎�����	��0��'��PN�}�e�nxBk���29���Ė������o�SH�++������N��E��aEĦW�Z-�sS_N4\,)��}��=J&��U�:f�RGE����q &��.�q��bZZ>�5�v���Y�!Q��V�t����M耢õ�� ;9�����E4�
�blY�~a����5Y��<VO��[�c۴!_���,��!�Mf]�-	<���7lM�T�O�67 �RU��)CrT�7{�1R�#r��B *�����d�:��Ӓx�rv��A��x�n�����ܱ)�	'�V�$��*p�2B﵋;w[(�
�� h�g�d��篘��#���
~�X�Qp:����i�%N\n������]yꂥ�+���f��<!g	?��_\�*�_��8�~4Q��4#9���Ju橇-����>h�PI�Z�Xi��M/��"Z�]�0a��Z)WU�n^�?��|�k?�"����Ȍ8=������_��C�F"	��ڪ����~pLx�zu^Ҁ�ia��o��s�Y�,e�u��5_��FDc����h�2d�����b����U����'$$��]��De�wi�A'��a	���,W�UGZ
]�� l�@q��[���H�6�j�]sEkUS��Y��*2,��a.W%�����}W�0=}��:*����P�EN����y]���r���an��K&��DG����zZ��uſ� 7V���+��k�q��a��&��l&��,rw�\�e�?��?e�-KDe�r	0v/�ey����ݩp&��+T��K
��	��>��<
��� Z/�����:t`^�!�c'v���+��a��Z�����a"���g�T�
A+���5�U��� 3�;���ȗ�]yz�+D`Հ�|��{�l�1J 7�����U-�hgH;60�\s=�ͫ�o�Ǝ7X�39�},M+��P������E������ڛ�6����K�a��J��+����]��a#�/�ve�@�X�R�%�v�����K�L���^�I�����f"f�?��Z�1�M��sHc�>X��w~7� �������Y^�,]�:���0$�ɋk�K���<셦U��U���r������k�ʉU�O�ʕ��y�tT���F��O��}s�ln���駖�}����Y�n����\a���L��7��\��(��������xC"�ߜ����	��2ߚ.f����S_֍�s\<����\|�� ��s��(	l���8u=�No��wb����T����D�Vk�[P�sMm���9��v&�� r�}��N���H��%_Q^��x�H��$�r�|� |�j���4 7���'��P�ng�e�<0�m��;�$л _+J��t�=z{G�r%�W}�h�5=�~�v�:�Q0�t���چ�2>��|	y��'�ז� �xd<1��^Gf��㺟zT��ps΋���4�]�[�F�$/�t��Yk�Yn2zp�������ad��/�n�~���S�NKƬ�zz#7��d���
�O��1��b��,ru�H�	�����Lb@��-�8fZwK��Z����7����䥝�F/�cW�%i�ZP9�O���'��dV<2�v`ș�e�a�@hC�qX�U*+�Ž�� T�U�����=����fM[m�G����r�:w,{r�yM8�N&>5E �$�ڡ�Tף������0��mVQ��:�@J�af��碑��<]��c��S�I�zCe�W�^��^bl��E�*-n��66���0�w>�iS�����n�O�2�l�ܬ�����jQ�f��3�T�i�A�cD|�,��AWx#���t#��r`�I�b�w[`4�;��J��������KG�(&6Z���f�c８i�K�#Lؕ
~$ ��i�wa��ûK? ˑ.h��5r�T�# �h�nF�s�2\EUG]_�ү��������^a::�U֛G�v��;�#b-�ӑl�n1q.�ހ�]°1�۝=�Ym|�J���B��!���A�$ک�~������ݾ6��K{4Ӥv���4\nE��9��1���-}JV�!�H���0�b>=v3u"�[�DU9��G����߭�k:�^�G���e�
�U~��0�b~Zn�?}-����:.�32�,i�	�F����������+�-��� 3�m�e�R�>+A~�'IL�X 4OL��!Y������/%��]���3+b����TS����&S4G�]ec��E�$�6Ǭ`�<��6l�+����Y�ܺ���u�D=>��3��G@�����\�� ntc���9����K!D+lp{�M.�Bd�ڕT��]��CƼ��e�x�������4�n��PZ��*�JZ(�T�X��U��LF���[Qn��noo����a��Ҍ�әO\~7������\:w���~$�9-�)n���b.2A�U��i�6����~\x�dJX|��h�����O��r�xC�p�m�`4�g����;W0�G�֮2����}}��㉭�� ݅#7�  ����$�;YR�y��ҫ���Q5��oH�C����R�z�J� ��"A��5�o
�9�� �kk�@'ehఠMh��������=�@�����eU�~}�۪�h��z�y�X��G��U5뷭O@����~�����,�c��s��k��/����
��/�c�i(��
pPWR����zMO�:] iOw,�ۣ!�ܱ�.K���k�A�ځg9�J4ɋ�*�?C�	��c�g��:��6��(XE&���8l~@�!gF� c.S�o�_>|BU3w�w��k�9�(ɡ��*X\�)5�� 6��ѩ�#JJJ05����>}�"��.���0KW;��-�Gm,� S�-{�Hi��~��ӑ� �h��*J��|��,+��+�B��z��q�?�g7n\·0L�?5����-��=�p�}v�m%��7����~u:Z��J,��)�w���eAN�-�x���[�+DFGGZ���埍�һ8����n�{�}����t��S����|�=@�i����K�v�4������-�k�h�.���%�ɽ�}G]��J3��4 �-�g��5!f����v/�i�@> 7�E����e�vs��!6�?���s?x�,�W�}(D]�d|��@���nȭ�ʹ��\I�($LR�z�3��
�q��D欿��23�J�`���ڡ?%<��H�d��6�i� �r�*a��o�*.U@j�� R S�(���%�FC��a��Csꦰ�G���4fOXp��xl�~�K���3�K\��<� �Y�ʖ,�:�ƶ%����u%?�z�Ԏ�]'�@�P�!}]3)��ߩH�s�kcAY���<��	L$f:qqu
��F��3��_K��-$;�3�"w�����~oP����^� y6��ϲ|>)5�}����nʚ@�(���+��pF�D-#�]Ẋa��,r"�"Y,��I�0G�����%���ՃmHy�n)�i�G�l;@6�-�(��(�n����X���#n<O<&%U�=�RX0��ǄΠ��2 gU��&畠h�u{ �˖����2���Jl�Y��̘L=tK�	���C���w�6�&w������U!�z�_�??x?v�Q�>*L±�6�X�	�yuE�;%1����G��&6h.m�����#���P��uF��lm���h-�=Wr��dZ�l��(��HN�)��9	-WçW�P+��Z�n'+�8�)�:u�Ss-�S�G�J\�w�7�K��nў��s%�Œ�����Ɍ��~�7n21�^_��3�N|��炃��e�Lԝ��hz'd1?�gØ����G��'�>;�([�&6���]_ǔl���$���םb)#���$�~iYvy'�����0mĲ^��K�(u��������Hi���)�T ӇP�X3�X�^��'w5��G�y��r��e|��qg�0j�(w9Y�+�0���c���z�U9�{�E!V!Й�Y,�`w��j����O:4��1\e�� ���9�&[��4�vxt��)#X��;N���0a��
�� ��]s	)|����c�
�#ŀ����9j7���R\\tH�@���"Wҹf�|w�0 ��l���+��v]v��V�Q.al�W�<]g��G�ɇ��7�� hRqw(�$��� ���$'7䩲n��s360��H�?�u���k�30�aW�x$�~C-�8bwʽ�(�a�ފ�1���7�h@V�,�0Z���PpGs��,��Z)22(B]fg|ް2�`���V���ќ��C��t��h���Xb��d�p�� A~���_]�줫��b���`�@g���4l7�of���rD�h;�#���������Hӏ��zu�aY���P���~0;]d����&�~�):��{tA�8��^��oa}Nwd6��,{�s̮
�Ж96>k`{D����S�w�'W�|2�+���Pa]t0�)��ˢh�+3�[@�-���J�@�-(�i\܇�R��5��[P5{b�vLb�dx�����3������6/��֧Y~Ű���o��<�ϸ�s���?�6�����d;�Z�V>l��;��2 �h�Q_�mbF�@y�;�o/	�n/��"��|w���1��N�+� �GN`���9�?�G��uc�N�2��S��W(���`َ���`�q���{٥Y$�I��< ����۳,�6�|q��Z9.�B�y���/ѻ�}��r����,���ᝉ�<� ���aN�oO�E�=N=- 5�)'�ey���<K�(��r⇛=LX�{����^�l���j�V�Wy��Z ���N��^|¼t��Z�tD#ٽ���������En��f!%�O]��$c��H�@�D��I�_t�f��ᆽ�$\Bá��ʀ�It]s��ܼ�z����A�s���	,�sP[z�H�Q�m�g��}u���$�@9a�OxZBv�މ�p�����bBa��J%iE�(i���F�8al���a
1����%�zxw,�7ғ�N�!�F��5u����O,����h�^5��r,'��1�\>/��+S�3�mS揞��"B�#��2�-��י*�,};/��M�h&,ՕW
T�W�f��+,i��X|��Ny�PAy����\Ш�MY���|���X~khl����o.4H�mF'���=�u��Z1���πK�V!LeiX؈yE��!F���p�8�mX���[�W%��Gq:��m�)R�m%tB��>��W�ͻ�,����n�z��%��U�e��SɌ�а�쇥M�h�x�v"ʶ���ڤp��Ao�9??lb���,�|&;�#ް�J|�i=�}�i��	�7?G?Բ)9����X�3WU���1��q5g�d��� &���?t�G��?�֫W
vG�r�DM���<)���|3�, �%�46d*�_-
�p��J��2=�b�} #�� ��2�YGC���y�/N�0Gh^�@��<�4+�<�7�]O����Ϗ��mJ=�WWXCM��1W����fF/$T�"�����S��7x��bZ0��m��%jjN������+K�r��X��Ht�&�,d ��9����g���q<1ȇ�X��pȋ�����J���_>�(Y1���?>C�:M�7����jqiIM��y�������ӧM`�Y*Mt� ��a[ꡚ���]���u��G�>�"���ϐ�RRRX����t�40��5���15eX��KSSS|=�N��i"������n�;3S��8y`ķ���أ�� ���5�4��n5ӹ���_�����ٳg��l�:2������S6=����Z�za��vz|DD|*�:����S�:����K.�@�� ���[�>�������J��ƍPu�:������:������?I�.ZR�`�UG��.�R���~�q/�g�Mx�`N�L ����y�u@ ��@RV?���l�׬��g�bb�	f�v��E�K\э������3VL�:��~����b�VC������!�İ�Ț�z`�4�����z�,��4�!|~�:�����K�����6�x9c�����bN���~:FM�+��kk�D`����[�/2K����M����©{䔎ԅ'�G�q��jWhd��Em��`]C֧i���f�����!XX%�*T]P��ǿ�t�����w��8�^.�Y0r��/|�;<b�o1ٍ��j{����B����sB���j�g�ɮ��n��p
/���t��yPHy��=�ɯ�Ŝ�:}����o�pW�g���l����X��eo �&�����K&I-�ŕ۞[8Z3Ʈ�P��)ϧd$E�!�2!d�0|����M�����1�1?N�h�:u�c��!Ë4�={��'��}j����w�+����ZX<S�k����Hj4�����9�_��O��������8���{<]�H��p1gVhu���M�gB��F��=�-��M	�N���>�4b8�������/�.���7�f��_�`aN�U��i�Z�c5z=�t��!�u�bX�g)�\/�b]���l�\/�#��
�u�2��.?�=@d��u�<�J�����~(o	�]����!jM+�B\wLmR���#���Ko�_b���vcR2��^��P��?����-����]�8�(��%��F�b��'�&�a��ȔY_��Q�QT����qXѷ2���#[j��+�m�U�aK��Iݤ�@XG+�2D�?����"�ǔ6y�P�;>�>�e�q�ћs�#������z��Ϊ
�˘�-��+K����76�0�������5p���Oh)�~����S�AE9""RN|4Y�#����!�Va�LPm#ɍ&���ݱ��!�,�r�x��Ҫ�6�������~v��};6��d`R"�}b�\6��*�a\��O�������\;�����9u=�؃[n;�k�n��_�;849��V�����7�/��]o��γ h��G�cG�c��R�����5�2VK
T���;xMh�ph/q�����xF�,�ak������d�#FЫ5�����Ԟ͘c���qbw�DzZ5�v��k<�������.���\��9&�&@���ϾS�,j��g(�/��q��L`0/QO�&񣍻��S�(Et0(+����ȣ�q&z����~�`;h��̖*+�F����|�掤F�: }��i�x�Ğf��gi�Z9Br�u^S�{~K^�d���":״�-�ՖM�=/z��=����Sox�f�;ƙ��KD�|�&�
���s%f�f�a��h�҉�&_���nrm��?Oh����kg��8E��a���JgS����$���7�5��|�n�ۃF����tN��ċ����Y�p�~�\����1m̔(3��L6*�����_m�E(q�y�6�OT��lc5}\ kM�Sw�J�o��I4�o�#E�� w���w�E֎��w��d� �Eҏ�9�s�c��$F[�G�'�z��ŠE�g��3��9����X��ar\W(�I9���)�/��329���<�5E(FoL��'����Rp����b�nSw��a���Ԛ*q��w���/(,Q  �'��ߵ.�jK�(#.gj���:Sv��N�!{]q0J��w�����u��c���q{�`�e���N��byJ�\(;u��c(W����qE����9:��ތib�J��\�|՟9$tt����|驒��ѥK���ۨ`]�8�S�8�;[�;�g�є��:�(�,����B��T�nl���ұ�}�ٮ�{��J=f������/#��/C�����~c����(G�׽QCw�/�Q�in�Xɨ��h�i��!3��1�G����H��SR�#ם��z��&���&Oc3-?��)����q\�͗�h,��N׀2�4���B�L�����/�Ϫj��C�0���/cK��������\Y*�x��K��HG?>��zzh����ūV�P�b�y���[V��bg�4T	���: "���a��.�J�Z�a9$Rz���.#��<��>=�s�Z�n�i(��/,t��G�����w��r6���OX���f�ע;r$�9B۳x��`3YqԸ�Ui �)���?(;�/���62�.�G�������	Fꚛ��4�L�L�H���yN^�+V���og�d�k =$�h��z���M]U���T,(�&��O�?s!�<�>g��tȚ"2�o��'.�U�aaCL~��[߻�����0�6�q%jʔc}��≧���L
���G �QҜf)��ŷ�Jo�lԌ��i���.:DS�8�җ��\8,,���@'�:܉i��.��$��ѧ�����!*F�Ŗy�j��k�̈��TV�޳���c��+���ruԲ�s�<@1K��J&��>omz��R/����O^]gp[�>�<���e�����ܡ�8^j�ZN�y�xn��c���Ԡg��H�����X��~�qK�I��:U�w,�$,��'m͹����n~�'���\��7��Ὼ x��ɾmk%�S�y?�J�wN�[�z�MZo�;B����K��zA��狠�r���H�ִL����:c�B�7��Ew���*��S�^�wiI-}��HE������[.��x�_�?��j� x�_vM���Ϗ2�c���W�ڛ� p��Rc��������:!yU��Ax���K�Q�����yhP�jj������K`a*�{���
�t)ʺ�����\&��/��u�gqG9�S~� ��1	#�>�;�^����#.�L�F޷�L6�Չ����i`����.��@��6?�!�X1��P��5�{%t#3+3�N�gd��)����墜"�R
CB�W���3l����P�Ӳ��xmyQ~J�-�BǮO�<��s�y9���MK���k��������l���f~��ɇ|/�����˾��\k�1���'�w9�Ȥi)�u�h��%����r[:�G�c��aRt%�6��w��$�ܓ���q4E��5D.��*�8h[޼�� 4 h����ђLʋ������.�+�����[$��&og�PN)ޗ9lq��3��f�a���m���j�k���.!R<�`��g�M��ɼ��L*ng�-_LCX�שc�npL���{/���rc�km���zU����.����M��Dr��IO���:c�,�z8��}�c%[��m}ֵ䏶?��{p����+e<􃳂m�e���V�S'�-�PZ�3�%p���N��y��ژD�"s�ƹ ah���%�z3�~���X��t<J��gU�a������g��O)�ѫ��]�W��QuM8�l�����6���+n���zp3[��25�D�u�V���� <�i.q�m����Tf
h�d�z&�q�������Z�	��M�7��n��ϋF>��'8��[�����~�x�Xau ��/<34���J\nߊ��;����J�7w��ᴿ�à�u�GP���^�2�u�Q9Yّ����7 ���R�gMUy6���lL��Iq� ���Of~d#Sq,��=B��z��aw޼�'4����ڡ09�#�e�2w��u.d�v:�F��Ε.����Vy��0�Á۸{㍯��3d��5�%1��gv*ѳd�B�OA�mN��ǡy�:�Nɽ�%��.�Ƃ��O�˼P����Չ'�_[b&Q�6g�w���m2|yt��d;Y�1���ҁ+��ʠ ��g_��y�}��Qx�p�������9���qV[fɢP����(ܞSRw�W"�9�eE�Po���9'9����V��k`Z�����h��x����A˱}�����D���a�|��I\�����Q���6�>�>]]1|�uN
�k	����ѿ����  *t�!�L�ֽA)��Z�X���uPl�ס����!WV_HI`C���_�$N���������U���݉�4��Gh	ҷj	߇KЀ�p[eX��ߎc�׍�K�Nm�%,��TjBN���� Uee'x_��#?���'�X�Nf����n��>���+6�S�ί� �Ѓ�SlxJ ����-�����?��X��u��B�Dq�R����ӚQ�,��[$���,�,տ'�m (l�v�A�Ӣg���kJm�\�D��d��3�C��f�[�?���a���Z��W��H+�j��7�����f�����$�+�+���s��8��z�)���������9�';l�Q ^���%��4Yi�PY՛�� ǹ,x�;�<].*��1�𳔝��Ű���T�=��F�����̹��W~��u1L��L��J{�8�%9��p	Զ� �T�Ib�,��i�K���.�,���}f#� ��j�f5���ؘ������	�4�Yei2�=���N�_��[V�(Z���b諙Ug7��J��lE2dh�[̈Ғ:uF���	Alt#ot���9�Pq���M�3c��b�G&4~W~�3?D��P7�1?����M���ǯ����9Z�t�J�S�9ӌ�]��' ����� NFZ�!�Â_K�P��:MϨ�2����0Q�XRX�,*,Ļ�ϫv�CK2a�����.����Ȩ:���	��[�~Z�~���Ӵ)uНB��ܼw'W;V�l���N���2�S������T�{y]Y(]���2�r��7{�}�(�3�TK&������ �$ZZFfl�2�O�0[>ۯ�w����FZ��ӋL���4:�����Wz ���U���hr��B�ׅ��N�'+k���0;5�¨��!�e�_�0�&�c�@Э]�_-4�F)~��@��bJū�U��|�L1|��%o��rA��ae�H��k}��gs�9��K�E����{k+��oNC���L�tD �%����8]�:�?���mr��V=hes���%H�N�ܜP�x�`�J-�O :��44}C�7��
Z�f�Ų�H3��fծֽ���HyI[/�ٲ��t޸���>0O{|�6AKYd(���K�@5��j�ң%{�O���](�6.LC�,��z`��R�U�Bsfa[�Q��EeMk�iO���!�$����7����|�A�z��z��ͫ�\��-\�����:Lf�8l�����H.�}ć4480�B�e5�f�ori�z�TA7��ɾ/�f�Z"���j���U�5q�C�P̡o#�u	(e'��ߣM|��m/ޯ$���S�ݠNܞ��Po�r�����TDc���ω\���V2��i����[K��v60�|�M���e<��g�6��գ3n�	]9ȋ�B�譧B���4>Ḋڀ�;Hç>��V�Z<�p{2�xptxГ�`k㫢J��~O��Zd�X�l���GpH�~��6T��
F=_HP�q�ؘ=;#|�Ժ�� X��
�KͶ���H�"��d/S̅L6��¯���Um˚��BS�n9�`���Y��RtPl����yM(�x_"����� ��ǤQ޾���RJ�	�8�zLo������'��&�Ͽ�Okj�p1.���������!���$m�P��kQk�!p�rhY�/���做�Y�E�lV364�3�%�$RM��]9��>���Wl�ayh[L�D|���b@����/#�z^F��.5�D�E�@�^LwC<����~	Ջo�STu����O_�Z�y\��ҭ ����r�d�TPAiOtQa�d,�u����ox8��҅J<;�7���	��BmG7rB�>q�3x'�#?��VW��uS�}S�7�q}�"^�o�����h�j*K͋�7��N>����`��jB:r*�Iގ�t�Xޒ�ox=���W�dT��/E4Y��JK�g����cCIiE�V0V��'`��z٣t� �;Y=��E�{���%326�j��w�&����:A��s�c��B�v.�`/�~.������>3ut��(آ^-�����"{5���O�k�߈ S�SGcq�P�����Õ��-�m{⃱� O,r��}f0/0��a� ۈ�^edn��+/JA���)�q��c=�8v�N��DXSS�DE	�������_)v��z�mo�����4��('�iQ��kz��� ��C���s�LE���r���br0�JuC��\{@���~;S�<����#kkkP��I+Q��vg�&�,���8�U���^Z9ʀ��]<"%��sGz�y�)�p���L�37�㔇j�#��j�"� `f�s��~Nr�}�(�����9υ��ܞA��ɩ� ;�e�P
m��,LQ.�����L���e�k�`=��\��cL�`�>��/O�G�_�:,4�߲��U�A�w�{�J�Nqhct8|϶��e�����긕�W������$.�fI����T77ٌ�=[^���&2d���w7� �,�	T�C@5�w1�:��G73�p����6�<i�w��׵%�6{Sw�T��8RN��Y�Zd��w�i��$������_x�z��t�LZ��B�8�cSSM����4�TJ����R�΂Y�/�� ˮt�5������lU VJI� 3�?�Ҹ`�z�L�v�U1�X�Y.[*���:���Ϊ]=$;z��A(�Qd���>j��V�M\+B�!�q��3��'�����ka̺�<��.�`K��Xg��q���������in��kd6ʹ����"����v���o_��Ӭ�"6e�3w�+綒��$W�0e�bN�;tNh�n
j\�1����oؐ��PR��h���e:5��Ú+�БԞ������ϸ�����A����
4�� ��D~5�>����!`�w�ʕPVڷ�,���L�\��m�m�RK���ճ��fz}][f�\@�JqI!�.(~�$A���)�� �fS��SQ�f-�Ƽ B��bk74���}m���Fn���7۩�4�u�@�V��Ե׬��6�~�*���_�犏Ss�?�,_e
4i�Y��+�2��@-3%~�-l$T},��l8�r��I�^�=BU�:C�u��Smm.�w�瑱�/e��7yҿ�I\�t_�/LZ��p W�,�l�Q{�)�EP�N���x�%�c�����oF�n�[�%/��y+�'�,��p���(3N�l�_?:!{4vښ���i����kB�7�� ��̰�*#�n����@ܺ�0����o�O��bߊ���WĈ-�]�5M�#�6�Z��ݦ��#��'-�Պ�Vz�󣏫��L�\@��Jn�ϡ�Tt�F�wW���W�6 �_y} �[����B�x��� /�wpN}��f�(O@��5��s[ӯ�B��&���}xX�$���T�4#c����Ẽ'(���&0�,F�����1�@l��Q�Ԇ��`9)�Q�Y���57߯珤�Ov�>��Vj��K^��Zl��oV�&�)\�`���"l��ky�ܜ�$C�Ceޙ�^O�Ϯ �.\�).�t�=n' �F��	���s#
P�\s���M�#,6�� �O)·��ty�[���-%E��Iӗ=�����Z��g>��Â�^��8���r=ӆ�>B���,D�����3e�����.��8�V2��d�#s�S�1���u��ΰ�C͋����;�aCc�T� �!��
�M�=$��S��������R�ƋC��W�f���ke]��}��S��yn��5㉌��?%�&�(+���R^"z E������6��3�2�7�
�"����I���|ҕ��8��7�Ys�:s����:1�/���7-<gvO�v�� YD,�t�����W젉�/" �����a[e 5R�]�� ?��
��D���
k-�WG哃)�!_?ݣM.`~�=�e�<L+�Z�9��({�Uy�T/sOÌ�N�T��4���eA�(��x�FX����I�<��qr���/��y�`�j����xpa�A��۫�qX�"JK9:Q�+bذ���.3� ��4�E=��V���v��F�z�K�>��#�0�R�bt|���,!Ҭ+��7�1���.	�S�������C�]��g������FN�-_�1RpU��1��o�k��zg�y6ۇ�ֵ+�c��[���Y��0��rD�xT�Z~�67��A�D(�'�>?�t^}��l�����<����E&�XJ����I{�/#�֣jDr�,ذ׫>\���p:����H�J��-���7�� ����3IM��(����`�̬�J���r���{,��z��xp�����ΞQ9�)�WW�yi��Ƈgp����0��\�G�gb�ڵ�;���W��cۈx5c�~�v�}�lP�������qR�y�w��u������R'�:!�g���QVy�/�~ݬ8|��L]
~ɡ"�,��]����S�K�[�t��\��=�nm��3�F*�i�
\�{��j�A~�F�4D}�����:`�y���1�JA���=��7n��#2|�>��sk�?��N���DX��A>|u����;�F牡e�	wY2_ `���A1Yӟ3�G�/���'N	
�����k��x�MCꔕ��> �>}?q3
��~���h���zy]�d�~������G"�Jg�`b0������--,��;뤾�e8�C~*N<���addds�e�h�_F�g���z��?1�Dm:�  _ 8��ܡ��{��J�R�G&��a��*�=�i�!�^�M�%���3�8�,T���Ւ"�s�<�}qcC[ꬕfc
��J�&��R�G�Ŀn �:CX0�y���l��c߯�K��X�X.�&��"O#2��G�%?��Ӗ�����57O��~�|T���F��7�G�Ё��%�~{^܀����ڨ<���-0kXJ�O5�M��u\m�۬���|%��b���:9d/P��X�p�� k�2� 8?X�M��3��L����&�ik��R�����Wןؓ��<N�3�B7�ϯ��x���<d�Թ \uY
t*��<�"�-�-a/StY��n|Xn�G�d�����+�{}}�7A�y5�x�Y]�|�,m	��>Z���/x�%�䤻O�s	�ܳ��ǍٱXR��V�y���U�����P�A鼦���5�����Q,oN��W����_�<���<�������@���i����g���Wn]��_:OU{�o����ЫH����
�*�.\�iiQR��n��6 � �ݡHw�t�t�Hwljҹ�t����Ͻ��9�Q���ff�����Y3�1<,?�L���b��Y����8_		���y����|�i��V	c�n=������2�$��ݹ���{�;�0�J���u�� G��[�������o�!@ۯX�gm�H%�(>�_=�!�?M ��-a�k��⇴��Q��������,�p��N��������f>ϓ�4E"Z�4Xy��¯�ޞ(������N�{���W�O��7��3��<z��G�ׁ�M%������\�$���[@*��惺�L~&h��V���~��dɀ���ٙ���������z�iN�e |c�q~<���6]gg���ݹ��0k��d�W�v���ᰝu?P���,/��:dI�~��_�`���6��i�����ʊ�u��E����"�ճ1"�y��G%M�'����ɘ�2oY���7�ܞ�9
1��������PP��h����4I-h?��w��ɜ�W��QiW7D�/8������~�T��H��㜳r��ؓi��F��`���k}0�Z5���r.	���, �B5@Ā���1��m<���	F�L��3�j'�������68O��
�"��{�o�W��i�J�TT:���2�ʘ���223�s��D�� �������G��̬��JDXXUUug��墽4;l#eEH��{${
i*��4�Qc�j��2(�}���jf�'�?jns6�`�.o�Eۗ�3ȫ������V�����{�Ez��1�����cBl&�CF4a�� =�,	ͮ(\��e���YG��͡�.�0G��ݭ���r�� �:��]5����o���gb+�;��L���7A�&ݹ��ʿW!}�j�x	2�;:aҐ"��7��'���Wu���T;�-�ȽO�_	�lL%�a,��FW*4#O5�v���le��f3�#`���~W��.�����s���?t�V	��]�`LŻ�+��R� m���O�l�%"X��؛��¦�; ՟�4�p�.�tv�F�p����)�K��W�Ky�c�k���I�������x�bzh�5�g� ~��m����`�?�E~�а�^�\��ՑV|go�l�>A5�<��#�c��i6<��n$��� ���0�mI�f'�=RO> j�;0.#�褙�G�ytAr�-L�]7��,��[C��0}�A�21,��׋̃�R[uͼ,�O�D��9�6�@��o��+}�H��x�({ܜ��U�f1|�W� s��$A����o�Bery�~��(c�*�a&�ru�0H�8��/�;�|Z�G m��<���Gz�,<%�����/*�'���
l.���L���^���̼+w���w��o���?]�Z'��^�9�=��[��ͷ����h?��~��C����H���xϳ���쌘�g���� �H����B��~�ׄ���7�f�7�$��͝�������5#��^zw��D�7����J2���A��b
�]g�����n�ܯB�bJNV��[��{]֤o9�F�{��Z!�"MMb�d�*�KR�˴=5��OB;k��8z�����[�]����t:�o;�%>��σJͅ���-f�����ۑ���̃MT��|�:�D�#P)�����,�3p����������`��	��2��^������v�9/�:�O�6�v�c�mS�|��w'Ap�ٻ[���f��1������7�RbC4D��5u�Y��~Dϙ�����A�����yʲb�q}
�? Odf���Zq3�>]���݅���{-T�
/=��x���xWo��>�	|�f�Ҩ�9���J�����0:psi_y?����e]�5U����%��]򖋇��ޅ^��e;U�k����:�� ni1Th?������I	
�Z�0�B��d�X�Qx�W�<�:u"��zJ<0�f^�k)nu	"�r���Ei,���_�&A��B�l&p��)���'��/�^����:���.��e�j:���ϳ���vTm���,�:w�Dޕ���qy%�.�����m���D�:�2Y��ƅK���<oy���4�ʮ_�ԛ��HIU=r���ʌ'���Ϳ�����L��x�#�x�i7	�S���&�˖�?�I��C%���{��gG��B�DTlb>VE����?�ə�t��Y�<�����,��==�}��wwT�BF��h�?�S~~��8F���O?}Ԟ�3h�[�5���/3�o�O�Hۈuv�Uon�s�������B�(���Ud�'��Sl�#�E����J��C���P��?���{7rjZ���\o�Ѥ����lh`k�,6a��"�c�k��h���&�o�����]U�W!6Dō��\}\s]�.E� �p�g��x���bn`��S�;��_������!?�Z+y����pv��t�<���٫B�\�+��Qׅ����D�;IU�MV�WOX�m�;��?w>���Ru�0�����,*�;2��~��ŦB�8Ϡ^���I�>γ{{ԣ��9��a=`8U^�d����������6[?p�X�f�dQ��%PeG>E���{2�z亢v�y徲�����j?[��4�y�A��h[Θ,+͈c����ԏ�Wl�.�������X�)d��K���a?��Ro5�"��A\��?j���\\HLn���l~ߧ�Y]����w���射شVV�%e��_W��_���Y�okwTR���=O��־ۼ���������>����Ɣ��ۦ�O�P�$��Z��j�\~NxH�6c�v��B?�W��@�!����yxe�����i��?��b�di&������p��4�q.�)��^��ﬠsAye���-�o������Ud޵�Zہ���	��)��*&4��H����`�eF$þr5{p~wY~�-��+�M�.����r�?	��������\�s[BR������؟.�P^�|�3W���� �E�}��r�����~+�����*'���ҒO��m_�?��N�nԦ�sA�c֦��W@BJ���c�7�t]cs�VI�w���C�Gū�24��U�H%��>~^&���u��,���}�(���\�������Ib��# �-�7��c�z���+�|�Pez��J��H��������� ^�F������?���
�s+���}ί>㏁7�G���J��d���D�g�&*�J�9Ѣ8��c�t=��xK���3:`�&0̴�������L:�_��r�*�.���nT�<�!���n�s��1`Se�����J�SK�R4�?z�"�ǅI����b�<y�9g�`Ҭ���&� x�E,fc��\���ޤ'���f��B&�h$�ҵP����4�#�bY�#�9���&w#FYJF<�cLLL�vI��m��K�=���#\�s�[;��ô[M12��\�����E�.�f�Sֿ@���m'f|Gܜ�c�Ȭ�lD�ᄛ�Iz�>w�C��SK��6��r2z�ޡl��VVRd!�\@���D!�����b�.�	�h6 qLG2D�9xzk�]�Mz���_�C f�ɕ�&�/�'���LMMov�Rds�R� vqs�RZ]��M�Zdx�d�>����`�|}����Q¿l �yJ.�0������ؑ�˃^m��=�^�ӥ&L�z�æ�f��u�d��bI�j�YcD�h�u|�X�{�|G�B�tt�<�3\7g����î�ꮭ��5�PPX(����o�GB�Nj����H�߰�Q�g
��;@�,Z�hB�fL��b�Re"��g��x�%\�;��!�H��{{t]g?�����+�~Um�T2go[�d6V�@o� ��d���9B,�y��i��t67�����'"N~��������>��+�ćJ}W�M�u�D庛<�����h;�|�A?~)��ߘ��Q��:���2���<�ӷ$��GTt��c�\7�)��$�R1(�@�P��ED|�:ْr��D�M�*|32(��`M��̃�&$*{�A����O���_���#n�����`d:�v�7_K\e� �����=�'��\Ć�Hg�Ҙ�?����qq���5�ۂ�L0�C�K�e�kͼ7C�v��q11��0v�c���?8O��0X�ЉY��f����O��c����i�B�I˳3A��4�ɵ��9?�+�Ǿ�\�͓&)l�<	qA�C��Z�l����j�z���{c ²���\}�WOǗ�k,�+�n��vg?�X�
 |Bge���_(�ԛs�{�er���Vh1XH[v	h����,@��\�$گث��QTV�F%wX�P��)&X����P�)1��Ff���iH߱s���R���O�U�&�YD�f>�)fc��l���b�����r��{H\�0!��ͨF���\Gui��r�����еD�@��B��U�R�lR���q��"v���Ւҟ!d�O�T�����C��^�r��{�6\E����M�.u 	��� ��zY9&��X��ǧB�g�����=�IIU֋�H���9�14k�-kxJ&I������q�͍b��x���a�>�����Pm�]����ށ��7�n����P��S��=/O,ۻ��Uڅ���U��ed�\�RVP���+���Vm�|n8mޙ&��ԑ�Q~R����M��B3��_f�<e�^{׮�a���_(d�DK"cM���Kz��}'��l�\�M���p)��j����tYf-9"_��L�z]��B��j�CǪ&�_u�9�q���y^By�,ߕ���VZ���$��g?��џrW�O��{zF��_�2�8��7��[�����5d��=չ��'��PJ�͞���.i�w����EMD��	���/��EE�;�g�i���'�*���}<]�j���� �͘&1������x���=}��i�+{�F�\��1��L:5p|��k�}JZ�>��}w��������k՘�r�9!K�w�4���C\�Z�l�/��3��m�!��+*¬hmm�K1�������\�?�X�/��Q��~	G���r!�'	$���`���?�v���WD1��g�o2����U�|F��@��Vo��S����TS��Dn� w>��T�!��ra��?J�V�,F��X�iS�;�6c`-��H4�H܂��q�`b-E��_��J�Ia?������K:df��L~_J�.v0��>�H�� 2��%9��Jv�Im~>1�z�z̻����N%9�l����b��T�������u��9�!@�7��Pe�c����-�{u�p��=z�z	�^�L�]�ۍQ�x}h�Q�~m�]yN��-&v<<<�J�'�'6�/_J�,x6 �	�"��������.��G�?�`�!�L�����#
V%P��:���N��]&`�74��7!Uh�ȄVue��ȣgc�'��̎��E�l��T�������.�K�d�<H��4�k�Ӊ���C����D�4mֆ��b�;�{�z$q�E���`FQG�W�P14���vܚ�?�ǟ��"�Am0_�.1�v�@���^J��e .2C侥~?���l����)��6Zi�����5Y�`(�6������Z��i{h����w�j���`y�����y���a: R+�ٗp먙o��;W�k��褆K�[F��5����������L����O����3�������rr�d��:1C�����9��b �I�6�oT#в���~����.�\����w�5T�-K�ģlR���P�ЩƂ�6ά_��$��[	3qfy��d?K?	�����-ֻ������gQ�1y�&˦c�i�e'Z����f��>%��i+#赢U�V��_�T��Ts�S^�0e
v����Rf� �6�o�/��L�������'azk��ܖ�<�"�	���O��1�[ؙ�p�6�K ՗��I�#� ����i��Ԩڭ�O��z�~�~D&�L���Xj]�m��5�VY,�W'c��P�;;LEk�8�G,.g*l�6����4hYA�gh��)�M��EԑkȜ�4�!6"i0���^��}�6����R�[U�1����,L �x��c|�J,�
�������edl,�|{y�A���M���X��~���:M'z�V���6�=�mwf)�,~)�]溧mUUr����=b����H@�CN�ό;j��	�gP��*Z?vu�� � S��5Cc�"���@R�U�����[10���X|�	�R �'
x5�`���D{p�~��������Jܻ� ���������XO[��C(Z�ﾁ�H��a�)Wy���Ӌ�!Zh���{ۛ7����wn����xnJ�Qұ����=��8��9��f6�x<y�W6W��k��D �6��6s�,%������2��_>_J|��:�@�	�(��I�V��}�K�"�z8��K�%[� ��Y+��:��;a��ԙ�<�
�3��9��:�[��kL����uvU��e����v��(��)���,�X6�8�maR��ׯ%��Z���>_��q=��4c)"�I�ߍ{J�Bh�ˏ*�&���աI��#�;���/�l)�4�f�q���a�`>�T���s�f�G���q:<2�X�x�V��#�f�X{:�v�/p�Vy���� �Pb���wJ��Z�� ���&X��������;�_t|҄�q�g��:���'[X��$i'�
N��~��:�N��i�'����bmO���)�ܬ+,j%U3;���Y��g7�6��ҭ�z�uבR�?�^}ͬ��خ��Tc��q��.��ָ�Z]_߾��Ml��S���� J�=����B�n���*������|&�N}$�-�=���ż5j3v�pzJd�++Y!�<�r/�ED8gyO�E8s���ԗ����]�eU�O��6�>w0.���ƭI{ �'�����w�[����~��M--�-<L`M��n�� ��<�C����a�(.;�9�jk�u�U����c�`�z�K|�iD茀�Ӎ��k��wu��I��S����0ԥd��i)�����q�$dt�o�0�b�;}��+'R�M���%@�.�YY��3ɹ;��DZ���j�$�4��n�H�y�<>H��ZN)�s��&���4@8;)m{�bp�YG_�X�#U#2T:��*'jfn`_�9TRaH�9O.=��S�虒jb,�ͤ�'�`�,��'~Y;�m a���o�<)�6���TΚ�[��5:��Җ�a7S�K"""�<�<���ɹ�_i<B���Om�.T�.(,Q��Z�@߷��>$��^Li�s%I-ʅ[eHs5���Fۨ:�y`�&�*q�jWp=�T>ބ(�۠��6A�)�i�a^�F,g���Y�������}좊��m|����\u'NQ��Z̖W#�nRn3��Z%�AQBBBq�е�~�ǣ*Sp販'j�lR:�3��j^-�'cl���ۥ-�t�)'��[�U�F9']�^E���oo�'����w�����
����(3���U�aw����<�X�&�N���z�r��=�0U�1I�u�2Y�r��$�;��aqf�W[(��L��s���U�ˮ�ު�X�Z�?є�/l�;��kV\b"��Xb�J�Q-T-��u���$���Sb5��U��V�Uz^��ݜ-�i�������ŏ�31RRR��%��Q�Ԋ8����g��jGEyE�����;Tŀ�Ȗ���t�ȿ������Ww����Xu�'�(�y<y�0������p˺�G��=�Ec �M�'�W%��+��s�Q&+'�Q���%r�j��m!��3,m�Y�j�;~��=�AI�(���"4�쏸[ �c0X�J���l	�0[7��kO-��ץ �����7�#�@t�w����ڴT�YN^�:�J�t\Ϥ��՟-L>��-����X�4U{c:gJ�_?���тMq�y1�����Ɖ��e����������O��6�blIy�v8	i~D�y�դ�|��ж�a��WCJg�׿
qU� ](�/:��}��o�¥oP��f�����bp�HP${����<����N3�1x��j�˛Ǌk��ܗ�g���fK���2>�� �Z(�M���3��n-����Č�j����`ʁ��|K�|[�j��P�n�Hu	��$ƺ&1�#�z<�xf(��#!���'y�S�w��5�#q}+��_p'8pG-��2�l̎UJ�?7��r�[�^���Ț�3��l�#
5)� ��jC%Ϛ�l:�}ijj:겞b�{���ǉA�[�s���RUEŌ��z)�� !n�+ϖ�MG�Sߟ#9F��J;D(����.��.LU
����q���6y�f(��UJ�7�܈QV����~�b�)�+��捰�Z���#�ْ�g��?Ύۺ|�W[�	uy:�=�~[��l�Y��\���ư�&)q�p����g�M� 8�������)��X{�ms��o�e0�8c�r�E�a�H�����(,mV�?�>�HH��3�Vh�͇֗@Zk����E��S/"q���T�����kW�қr��cAQ@�ޞ㧰�}nv ��J����!m������Db�[��|�<�|:4�L��������h��wn[�%*Ė���Փ:�uS �$�q|�?h9��]zh�N��S�G%�+C�%3�)����>?���	�+"=�J�.m�q��y�F�a�k��;�����^?�{��<d��4�x'���}5[�{++|��X�8���}n�#>I�k3�"�4��  "G�nwA����9Q��{�+O��pJ�u��(�2��6�L���o�u�N����y889m�,�g"deh�?�����z|=������Q�qY�0�6J��J$@�aY��߆� �f��)��:��X<)읨2R�R��`�#���§����̓�����vֹ7����<�s;�d�\�p�!�O���pR���tOC��� F*�\�)���fc\ϯ=�cL�*�eA=!�/E˫��v�T����B%*M����Õ��IpiG̿�p�jٸ/:}s~*D�8p��q6�f��/J��e�3K\G�R\�VH��C�^�=�^�pm(vt~p�ۮ�E�gK�X�\ߤ�ء2s��W/Z�,���s�4'K�I(>TC�6�0�������9�6�Q�&��-���{t��F��7�|�_�?����[�z�n������̃��);��n{��������xM���VC���/�����a���=�����Out���AH��u	0(x�H�PM�pN����us��[������"`׃��|��q'���k����q���^��P(��Lk75���ݫx~O����~��ϳ[��U%1�3�9n��2�T��W�+k��wq/}$Q��]�H���h�DN������fv��	D��vhppb�c��^zOOǂ�Ҥ�WS�h͔p'B�e�ޗ���N)��aX�>G��e����k'><�Kj�����|?�U������e�-E��_��5�,�
+h���zs�_�T���a����Y��R�X�|�W	��W�o%���Y��xH~�K��n6oS�r;qx�c��ٰ11}�1t��P��XHH�5s4��uL�\�,�T��O�t�i��]��\��5�e�^m��6��ko�G�A|��.��tx�{{�N��p�>¹����\�NxX9u8��C�m�=��O-�v�"�<�<Ŷ<E���*,�B
���)����sDJa @�9�,��~1���l��|��+Vmr3͖�� 9qr�4q��tg�Þ�^h���X�����d����M9��A.1H�E�eU�����������*�׈A�u�B�Q3�H$�-�p0e��s� _�{�zo�]�}������uXU�k���V���ƭ{�H��Fr��MEbF�Y�����[d:w$���)��PB�!ő�����+o��WUʬ B�Y����8PUYO��ky5Ng�?i��8�����~��f�����������2�L�6�fffX�v5110�ݙ�Twp�kgY񀛭�)eZ���#%*���h��h	)Y��=wݦ�򦩳8-M���a���-�\�s��-��Ln+�BU��m9yz�(�]B��m��ֱ[͛�\��Ȍ}~�N�z����d.��K?B��K��&E��͐ok�a�
�6#�[Kr3�@�{��/?����6A�ynu��<�0�f䃒��v��r�9�ŧ���UM�������z1���,mT�O��#s�J�4�����V˶�j6�ѕ@����q��7<�����f�K�2%C_��밪ss��1���)֒�At�\�>7��@�e0��C7	�U�Y&��Y*H�/9B���B�v�	�-f�4,�:v%V��{����0��8;p~��C�*�T�]�i��@���g�+[~f+������`&ʅN��j�F�*���*���M��[&�����͋IBǔ�p�-Ug"S������w������d�̰K<P�6���E���,}Z�)� ���H�=9�[�ti�(�S��iy�U!�W3s���^L�:Lou��u	�H�T�vT�R�n�9-
h��ʇ�����pFH��~CܢPx�b����)+ҙ�H�ѡ�Q��H���*u�zSXi'7� I2��������3Q�\�,
i��X$�Y�Y�� ��1�Y$˹��B���Hդv�ӂ��-�:"wSs�L<8WTS���&�b/�0'P��/���%i�p$��| o�صXC���@Nq�#�%��J���R|p���3m/��4���e���<F�ߺ~>��U�"m^��+�E9BWg�?�N
���Y�֠���ܕf��}D��G�-g��|iX��8�bL E6A��FN_�m�J�� �{��4?�+��.��s����`!djB91+[h�*|NthߚE��3�P��fK`�h�X����]@�ި�z�O
L��yT��[B�K��&����WU��y��s��������2[��(JNT�N�;�g�ș�A'�rgV�.���ͼN�L�vؔ�G�ݬ���j�k ����)��-X�f-E=a�8����R���]���������\S�@ߢ�#�����<A:���Z[�>�ZI�/�+�u�T���>�OZ���<�r�$����v����3�h��:�+{W�S���	�bS	���r ��I���Ղ��.��첕�k?�w�:�>;��������Iܑ<��S�s���4r8��������|���x1��F��}�Di��L�W���#L���R���4ΰrX%��@*�<Nq,Lv�`�"�7`��Y�_[ѫօ��]نϗ�TRGi��;��o6��H���Y�!r�fMq��k�
�{�U�`�fA�!F��)l.�kaS�":�y�v��m.�||�2���0���-s�� �/�Fߐ�o�-T)Y"�[6ww�y�i6��\&rX�R>I�}֌	��M�>�h�ۀq���d��%���N�˞��ރ����֪�q`R��+E�.	D��q�@F� $�A{�D���q������i��-t�ZU����PPF��E���!o+2)0�-r�R(j6-�ۗ�>n��|���D3��À3:@S�Bq�2\rU�!m�] :55��������EW���ЬL0�E|��v���?6e�*�{������
�9g����=z+�S2%�\t9P�!�:���ou8K&QG��&[*E��:k@*�m�R-�d�f���4�hyt�]����D�TP��z���"y3�b���8�&smmn2󠏾GT_y��A�o��*��@؜�:��x���*�U���:/\sϗR�Oh=�P���mSs��$�tD1��G&����ZY�����_%H�*�B��h)����rC�^[��Ig��ӓx/f�=�XC��$�$(�*r<�pU�����e�QF��KF��W��e���@�����> S�]$tJc��d?2�u��u���|�\$�z�~RP�}/�Vs���
DC�J'�^׋kT����8AN��40�h6�ظ�Q��Zߓ��.�O���<�e���]�	��(�s��@�n\��kaGg<l����f'�u���r�D���b-I���Rf�C�7p"y��n'�~������Q��0�C����a�e��{?�k�4�g��ە��hn:�
�����{��.JA�dp��
�==8O��!ycc�U�/�Ү��q ���2Q|��U��7#�z���R�bql*	w����)�ө�߭���w�������^��?OTY�Rw��;mr��@����}�/5('�V�m�XF� ��l_��{J(6�H�;���Aj ��rRx���>gAM3�0&@Q�!?�D}>& �����s8z�r\f�xc
i�������?� ���<����&���!z��~ޗ�(�!�����~ǂ(K��{	|�����z8#����?0��1���8�]) �;>��(����a�I�@p�w��ưK�<�7C��f�� ���B�L���R8��UؕMܼ�y��!=�W6ujh��[��O��O0܀DUP�
}
!�,�Vm�Q2H�6���-�h�J+H����i6�?"�v���I�_k�J;�ڮ;t�jf�1>2!�c2|��J�y��K��Ιf��Y��)2�ҶA�!��F�*/��s��+A˂��'M���l���~�@�w��<H���qg��v�����F���T�w�#��Nn�x62���gO�׵����BU��Ft�v�m�����H�N�7��'qh�9�Ĭ��������r8��ZQl�u��E���8���0b���|kf��:/5�lđ?�X�(hЙ+y������`���:��|�1�:���א�`0t
D�տd�ʨr�!�D@J�^x�+,h�1�\Dev�W�'2:r��A��ߖ���N��94:88��[��b�Aߣ��x��x�X��ƣE28lE��
����\�]�AF��?��9��.U%�q/��@B�_݉���1�2/`|6�Ȃ�����]az����|	�N���	�W���{zy�N~#�=Y
oO��6��F��Nғg�M[O?���k@Y���ЬC������������|��qV/��4�P��#��(HY']>,^�.�GwkW��yq�#_�Z�GZo�_�\1��%�>_^�Ϧbh�R`^����ܚü&"��?��x*<��c�����vi��#�/����0�LVb�Y1ɚ ]eNNu��K�l
 R����
�Ո�����G�b�/Qa[�z�z�k�]C
g�*k��t�qga��X|��v�]H��" +g�u�����ɱ^2B�s"s��/n�P��m�!��3M�'	�d1��{�q�}�%����P���ԭ{��9�y�d�\Xyꛢ����`0=5'(ٌ�� +0�o��^(�b�Ht-B�o�<R�"K\�L��h�ɀ�|�HM�/�tߪK&��!������i^7.s.�)9ŏ�Q}c��4߬w���F<y�VV�k��O�$��˥���f�D�� �	�
��vX�F����[ϰ�qCDʂ-�J�;/c�Y�c�fJh���Iqw����m$��
*���
F�Y�����b�$�h���&QÇ�N��N�界'�;lIj��0�ӗ$X/_�t9��C��0T� D0f����)���C�f�F�*�{?ࠟ�S[ac����ԯ��2^����Z<÷�-��7��(�~͏�fz��!�A�s�+������p�Q�H#ݟ��Ujk*�Bkm�ry~��U��a���IV	���ң`�ܽ����2a#��V�}� ��~s1���W<5�[��,�@�C%��J���n��#vm�g��8t[�&��n�m�H��H r=�OuG�!1E��Ub�+���1+�l�m�	dp.]�9�-◒�{�M3�i�	�ǻv@�_�w��?�K�5>s�~�<��"�F*Ho;S���<���G���Ur��=�V�N��dK9���O�OC?�0������:�>��<�R���2|5I�����l�����#ۤ��ފ&�˕��x�M�����[���X+"Ф`����Ԁ����}g���0�#�����
<�>��k�k�ʍa�zH�9��I�����OQ��2)��
&��i���3�	,��?�a�� k�Y�C��B��$���d�-pRʓ���.�E��3� ���O��� ��a2:�M�z7e��Ca,�Oo	���d�l�B0�����-��j�.���nT�>i8��VEt=���<���P�I}z�I�_��/.��N�.��u��x�ÔaLR��D=��-��W��pRӱ��e��(;��+��	�`[��� \XB�;����Q��+q�ۿ�q|՟y�W��͆d�&T{5�P"�[)W�;.����&��ʅ�RXFL_�ig�?��@H���[1o�#�������?8���`��GD5�[��ζ��v��6����X-Og^61* E���4)�7��:�]"��_���<�ev]gUJ����U�r@���p��+&H�IB�e����"�O�#��?v�P	���h�O�W#)t*�n���<x��B˕6�؁�>NiW���'w������v	�|�7���"R�~nxd����9���~���)Hh�"?Z�n*��*3�N�j(vb���ټ��t����{�.��F���i�`��HF��|-�b�.��J_6�Az�q�E���ZMڞ.#�Y�vD@��E�_2h�M���?dl��A�Lg{���C����B��-�h����>R8����r]���2/�+H_d{F�n$���@z���a5���0�������X}��̉�5�cp��m���ÿ�[��@��)ֶ�Y�)�G4�{mk
�ޛm�Dh,��Ij�

�JG}�/Q!>��o�����|����!�D4�2����v��|�8s�K�'�C@�O�E�i��@<� dQ1'v!x�$�RknZ�0NS�)�:=T	|͍�`b������}Ľ���ZzI���)Z�F��w�IrXd�]�Z�C��q���A,�cG<��!��{ܣ�*T.����%W	bͦԨ �et �B���r��-�j}�:��c]	높�@·F�o��Q"�d�����{�?��;(���1Tك<N's%G�g�1�#��l���ޣ��^��r���TY�h�/<���KI��2����L5ͷ�����@4,H;Ș�)��z�-Qh���zU�8Z�M�_=u�E��T~�faY1���V��uj�J�[qg��1�@�P�E��9�]Ƞ_|~G��*�v:�X-��Ǚ�P�R�����N�`�˗��,a�'	�\�6q1��|ɸ���C�R������"@�[���K�W������W�GL�f�Kq��O/�~ ��|��U���j��R�?�F�5?��0D&K>}��{g#��������#��@�� ~���LY����(�n�X�N��Ց��c>8�pHJ����dQ8[���e�b�~��0��qe��0f��y#}$��:r�}b�4H`28=<z�_?"�y�����t� s���ӓxq�p�+����&HiR��p�������c��ܛ����s/�l}�����f�Ar��ɼk=�Z��h�V�Ն
֦���0������.Yx�IN7������?�!�c�� ��A�)�-Wgs�\#@ �������������ݸ�@��NC��e ?���w�:�����"����"�sֻ�s�!ƙ����Z�x��<�{5%#�5Df�6�-6��ɾnW)m�޽/Ho=]x�
�҃
ec@$�f�xy<��, �g���p���8�W����<\C�p��L��#�qz�zJ�[�0�U�u�)c���뿃�u���7g���I�6�O Ja�?g*�A�& ܦ�����g�T�z/؄3KА�_F#~w�S�ҥ�����=;�_}��N~o�t1iyx4Q�&;b�|��i."H1V4������pʹ��P@��lQ��ޜ�gM�t޻z荧l���\��ԡ�I"݄U:����1���Ä�GHt�R�7�ܜ�9�n�`��˼�^FQ�kd!b��=K#KxR����?��<Щq��,��d��fPi?�7`�x?�%�NM%�b<:F�-���]F�8��T�yO9$���z��&���n�&�D��v���e}KO���F*��=�2��k4�(4M:��5��Dz��������Hi��.��`��<2b�������6	;����M��YI��r�z�p\���v���/:��nJ+�H�������HV�w"F���[cj�)p[��#*M>y�X�4�����%s�d�	]8b,��{��-��}}Nh�\��������Mƙp�����-���ň>�����·�Q�.��-��E�]cn�'8�"�#�ߧb߳��_Igcb�2��b�E�P/ffE�11ύ����������晩V�\*eæ8W@@0���q"����<ٰ2b�(�!U8� KƩN�Fy����bA�)��n|��ǰf�t�8�g���3�5���
����0�����m{-5T�Glrv�>�&��_��aVT�XH�h�b�Q��N�����Yܹ��b��c�A��@������3O��(T�
+������C�M.�(�2o�T�֎%\����#�k�݋cg�6��;�]�m��:�7�/b,A^��v�˘o��#�{~�lJ�hsN����!T�5[稳�wd^^X?�r�.��E s �rw&�cL�6��	�y��K�		y�����E;1�k��L�cL��gO������^��zQRZRQ�Tr�P�_�Qrtӗ�v�@��6n[�=1ꇒ���n�'�(4�� g�me�n�BMBއ��Ԏ�NB[_��_٤�_�jt��a9���{w��E^������k���-&��N}*�B�l�R��C���pG�_pc#	*���(ǐ�=d <�T+#�s��5Ӯ ���#2�!�������.$�}:N}﮶���~R&�ؗ�x��)�SQ����A\�,�W��z|&���l�4��5�� 2b�F�ܞ,����pOY���֖8c^ӧ�ɓѹdB��ʻ��1�7J��C[I�q|�֘�gc-\cI7��e�|�eY��R�`�����u�ch{|�*?��V�؍�<���E�骃��9�>�mys���F^�S`�=R�t�p.>@B���,�<ڃ�����9?$x�#��0{ٕ�?���ςB�4����LF֦��ѭ�TG�d��ۓ>����w���F�q3��kJ.�e$&v�N+͞���������١�f��Q23��l������D� �A�*(�Nif�o�o��eʣcl�HO&�o�zbI���H"''���j~�vp!���J���*_���W�x��ɓ�,Ջr�������Q��M$�;�Z��ʼ�"&vw�ƈdl�68������A����~ɬ_^�zZ�@�{�CO:(H�coe���.��ª(
(*�te���(�5t�(H7HRҡ(�� 1 ��H�P�yfpw����w}\�׺��<'���9�9Z>����ط'P�hO�{aV��"�ы8�},B��ٓ�B>{*]㊔C"YЪX &�-7"��T�y���Em��1p�N�㞜+~(F�*w##4yڕ� 鵲K&�����S�+ccoq��z_3�/w��<c�-�U���=HUQa��2t��� �א�S��/���o|�8j&G������2��>	{9�,??�P)1��N^&�?�8C��
=�l(iQ��������斍����VV�c%�{No��N��iky�<���� qs7k-*'�ɫf�A>�Q�[���'۠��-�»x8��&ڔ$S$a�\/���Ttx��ۃοǵL���-���*�lܙ���nuZ7�=�uzX��⣚��S���T��|�2j����fo�������-p4uߘw k�/�������E|��j0�s���'ߓ��y,V�6���\o��7���֛^�!7o�{�*_���kr�w쏫�A�G7w�����o~��vn޼��cF�Հ[C����W#�'�?�¶i/�@ޞ@��1P�2��ҧ��./���sY���[������J��?����9*�Nr�Tk	�f�)Jct�������'J �~D�,��g�/�c�f�L����.���s���BM1KΓ�:/p���x�)^� ^b{�ɠ��lT>$�pP�M{�y��Oѽ������ـ��o���$�� ��ވ�Å� lP�z8���&�Q3����H��*$�r�3�&6��5/9lO���Q���{�%tU�h�Y"C ���U�6�\M�����i�t���@V���߽�N�W��S{Mpy1
N��/�钒�v�גb�F���Y�_��_0��/��V��.��ʨ/��y����D���v���k�p;�X^Lm��X8R�����A[��-���TrJ;l����Fי��
��Ӓ	�+F�5��s�]��0Y߿��}�I>ȷ#�O��u�힄�¿X����	��~��M/C����M�ʇ5�ɍ��|�*�r��]�4%?_�E_��[2�p��3��v��89hk���Oá� ��ʶ��$^�E�*;G�8I����2 5{��y"V���a�Q�fn{fw��y%�������G��B�`�2LG/��������ך���e�Z�v����X�J�xO&]���FNשP�fJ��3�������%���qÌz�:,����[]M_�r�6��X��B��ĳ!�н(#��"�yV�d@2Y �񩎳ʥ΂g����&�&$ǭ�z���B�����M
�1�"�� _�e�k6������ߎ���z�^�7
�T�ۓ�o;p�x/a20y�v?3�_�l����͜���6^���{���@��f½>��"�?��ގ�(?��|�/����l�u��f�L$��b�ŵ���$����q���06e%�ld� �����������}�4[��N���S��ЫMg}�ɾW��n�]��/)�M!9�oL�f{�AE��l�z02�݁#���8�����O�H c+� ᑺ`m:B�\�e�F?� Mu�$�]�ɣ���T�9j�y�'3�2ǥZY"��i�k`S�
���� ��6Mx^{~N O�(cp�%r9�Y� �Uź�*:%[������ſ&���ń>������Իwn�^ݰF��CǱY�t;'�!s5�5���
�*��]�ܓl�/�#+���r|]'q<tJX�� ~��J�2��Ւ���|[�F�a�q@E�Β�wc�9���|�����@}Xν�s>Z��3�=)��k ���ƶ^�n0rr:}&��)�� �h��/�*0��?F�ɼ��z'Ɠ�F��nll�׽���E�6n��d;?G&�h��a�Ò��"��2�ۍ��(IsVJ�~�S���_e�*w�|Ww|�v����ER4=��҂��rE�~���ّ��]v�a�|��I�4^;��F����.�V�Xu_�̯�z��^��i�Ͱ�u�ō���J4 vjּ��]7�f�>\33H�ϊ�p�D�t��vh�43�Ȱ�@g>*��`u��L����뗁�Uq�	I��j��܁W���lͳe�,�(�2�0&��g�u�+g�� �~�|����&����A��0R�5��&_��\��JX.�*u)e�Y㦶k12�b�Ŕ����Hl�\֘8f�q�^7TY��@J9I[�k�hfd<[S�5��!]��`I���mTT����Iy��?���S�8*���9-3��!���X��^�f�1=
xr��oI��/{Uˤy�W��C�+�/������w����G�Ye6�2C�a�r�]yCQϷA��l'�$ϼT�Ҿ�\_T�닕X�S��հE��J$������ih�_��	��;��۷���o�{���d�UUq����6��wLw$���srN�O9]�h�>�6��c%�-��ځ�"��H&��&�9_0�crWt��Y)u���� ��2�ÏVL��,�hPX��Sl�W��̄���p���=C�7��_��1�nZVq���Ӱ�ͯ/��/����`0Y�V�.�`�j�d����Nb| �D��]0����@�\�;�I�����W��iғ�i&����u�/��G��:)�� \��Z���o<��d}WG��ܝ����Jy4N�����1A�/u%�7|��>��"���Ɵ�)p��prn���+�i\���X��w���rT�<x1�|��-���jW������9�;�gg����?��E�_�t�g!��D�f��|N������SM��&>�Q<����TmS��9��Y��ۣ=�1��R�,R�Jf(�A��C��bh@-���v'��{��n���:�M�H�0�s��'?��g4�mu�hi|�����F��{����v���n�l�	}����ۆ�2`҃���&�
C�Lb���6Dqs|=�_g�Ϫ,�wn�I+ʐ:��v��OM�o�UO��k2�&��s�?�{����d�J&�&�k��ܛh�禨N4��̎�Dr2p����mp�V�������B�t��&�wM���=1�I�E�8��כ�t[����� �<D�)c�Ppڙ>���0�� ,+8�]���/Ee�ѕ�(��H)�g!�9�e� �q� Ɏ��B�r}�ǅ��%����t��!Tj�z��BT����R	���O5b:~ֻ!��C�����;��^���:m~�K�\�3���-��Ϗ*����j.��I�X+(����8u�� ��r����dg:s�|ɛU=ޭik[��zQ��3 ����\��|cϪ�����Y��u�	aO�����BzgYIq�B�q�ݘ�T�~=��]xUM�\A��&�3�!���A��*��.6J�fS~�OU���&p?��?��`���6��J!��ԸV��k��+���ʻ庬�oT��٧�P��{C�+�c<���W[�����gP�-���/� ��FG�����2g%M�A���rKĞ�84;��0��~v��er��� �,����rMb 7��ȭ3�L�9�MZ��1-�`��
[B>ǃt�JH�.��b,*�˸X���%�2���/��������Ny�8�|v����y��əaY�l "sN��(�� � 9�������	�8�-<���,oB���Թ����l&ϖ�^:���ё����(ȎMw��w1y )�]�ۤ0���vO�v�B���q�*`��sS�b�mmѝ_(�~N��x}4�+	��?�]P}����2 4��T�ТU�����.s�K���C�ځ��񪂣ʴ��a��pQJ݋r��ni�gk�Fgg��L�ͣ�Z�Dy#�������Z���s�ˎ���(�����ݓ-<�a6 �A�c�w�FwO��Y�*�����v��E}+�V8�����e�2Gii4 e�����F�ltG�A�ri����H���8oC���-2N���#��ґ�Υ#Q��X"M�kjp��nvE9�k��o�F-������8�U�����!��T�"-����)�c�R���v�uȧ<��
�s��{�
�9u%%�sWzt�9Y˸�M<�(k�6�i�l�(���Ȑ�����L�SZ�o��X~��D�"�a���8X�ʺ�7�~���������/n�H{�"�ſ�N���9/ؚO
۪�Y�\*c�;�OO��� �Mh��y\���߽i8�pz�l'�>��'�H0mҕ�_s�:��t�0IOb������;ɉ�eRoj�㣏-�ǆ���K+$�n?����+�d���^��%_a��*���h-#��E���ץvG���O�@�a�H�=t���8�]Ü�L�g�AQ"`��RJ��Ʊ���d����&��B�/����O�����qո7,���D���S�A���w��Tsv����s�r�����]���N��*p8;3�����x�ˣ��I�uR�\ҘN���3�^�6q�o�k�ſT=Q��_��?aP\����[
����F@�Qu��8G̎!!Ɋ�׬�bd�+U���j~4с	Wc�|i;��Y��S�~<d�K�� QZ����"���0�̔Cw��4�����SY��*��2��s-B�=��o���BM�zj\���lUA�_7�R�W�NQ��An���m��c����+�������;$Fגb@�	 ��
���s���"o�7/S��ͨ�.>~A�-J �2��?���2ZQk��,����=�a���<�ߥ�N����-c�{��`=m�i�	�[���w/�� �OE�	 \MG/{��r7�/o��f���}���m������wc.ہ�(Y��{�Q�FF?^.��ܶrTp��ebb��P�W�s_⅑y�}�'�Hdd�!j����W� ~#g��ݩG*�?�=�h��˩�r����ş>�}�_�=V)_2�Ҋ\OOc)�p�����oo��ۘ����A���<��5G//;,���!Θh��Ң<�va�����WE��̣$oNjiiAۆ�ڸ�R���{���$k&�=\:r�	7����8<\�ҷ"XEmÜ6@�j�V�0�мx���3R4�I� �z�����f�w�7 �9�Y$�d>_�~
�������RhD7*�#��o�s��Q�)��� ����r{��R����S��:�}镙����mqW�`�l�6;���vA8HF�
뮤�!9.���H`�+]��G3;x�ڳS�Q��(���pn/�[q�e��ޤd>���Jqi*�I]L����L�(q����]lW�������'��A��_LbB|���.ALU� (ћ���j�!�1@'�K��5�BTT�X��������b	�T�*,�i_2}N�nV#�8��N0ɅY���`4���k|n�J>�=����w�\�S��.U[�dK1%9R�jeڡT��|sb�JbӾ/���=Z�����R�f;��eҁ�(�Bd�Ez0��o�,�r��t�Y_8ߊ���wn�
���"Y{��/����
"R�-�Av�6=G���,[7����K�=],������ ���0�5e8.oSy�ק?g4��F)\	�:����6	��;�>�S���W�V���V/���'�HInS ��~�|9JO_���W�)d�?���̓8��X�1A�z��P�8Z_6gQE�N9E3D.3@і���Gٓp�9ts\��$���Y�O���"Ɩa՚l�Fn%%*X~��|�1���{�;�;��n?�,Z�|�W�_��I�j�B�	�v�����+�*-�d*S� F�	��ε�`��w+�m��g���N���c0���em�^ةf�L,����E�.�IT�U&#��f������ў��ש�4b�
��(M�?K��Ą�g�N����͛7�o�q8�J�'f�yN�m�NN_t$Ԅ����M��f����(�<ds��j6���P�2[̔��"D�=oĥe� ��=C����_�����%���A��2����7Eoz}�>HKK����y�MOO#�I~�%�k���[uhM�!u[l0\��_;R��K����&��#Fs��;�!|�߇��v�<:V"�-�"����ڬK9ݭ�E襤���7r_)���d'�_�t��$���*��R<�y�a���������!d��fSㄺ�.DV�+Mm�Ob��<��F��@,�I��xl3{tt��P�4ta��Ȁ[]�++���2C��9v�UL�1#����y�7���K��r�z�����/�K�`m�<]@�@'?���Gf@
�Xm��$���h��(���ț
f�Y���o�ӯ��Yqqq*i��ڥ�Jw�u<��m�DfK%�}���NX�Z>+��y���z���ȃH��+Z����%R	��77'kkk#[[��q`}���$e~]]R��	����"����[�="Ĺp�?;�D�uu� ���뜔Eo����Ï�4�L�s�v������u�ذ [!����9E�C9���@q���\�vz��j
E*�w��GD"eq�W]�gL��o'˒li���"���f?�Ɨ�^~����5׼+V�.�ao�x��"�FP������b�طU�f�s%���(V��i$S4k�����?N���[�^�<׫��˯Xc�l�������oN��q"E�uڷt�|�^3'�@�W�!F/;�I��o��� ��!���.��f����iC-����&��6��:����G�����'�~t��o�E��]e�2wRoD���<Ue�鵘�x��+��V�]�X�g��J�{9��c���$�>G�P	��q.��7�?��u++�,����]��jy�0n�5�VKC�N�l�q�߀;���%�+���c����\g,Ȝ���Ny�y�g��b��(m0��*��2_SBv�?���a=�2�
������+Hi��!��,��-�3��oT�ް�}�iYW��]Wx#������|�H�e��Q%����_��K,�����h������>��9�Z��S��1a�(bbRK���=������L�aO��Fe³���Z���l���ݛ�)n���b=~+�9( �|G��6# �x��w��+e��]����$Χ8v��<�y�������H�TLL2���3����� ���~Kǲj]����������ݞ���>�(��F֣�6���W��Hi#����%�;��rP6��(��1=k�'ȉ�fޝ�Uf;{�@u��^�qM����a���	�I����@k�H����X[�'
؂�|���P�}�9�^�c~��*���Z�`��=��|����ƫ?�}�������u����܆�t�W�Ff������I���&��f9
��-K����0e#�9x���=�{�3�cb�����г��xO=��"�(Cjq�hL�R��+�P��a}6v��S�N*�yg���&uC�	~e)  N���I���#ᶳ�sN�t�e�!�n-��� *7�̈zu�6@�����s�"ʀ�z��P���,`ڀ���z���i�˺�&�xK+�Q͎0�o���'��A�}�@�$�o�0���G�*/dbFzP܀
�5��EE���2�|�z�x�'�%k�Kc�/a-�i{~o�x4�������J�;dpp�pJE��S*�~�r�	�a/����8k�/6l6Ҁ�Af�:E8���ޅ_��_�s�;z2ˍ���5� ��au�B��{@[`&.�y7��"�S����)T��Ǯ���j	'Z&x��L�]0t�A\g��SS�:�.���T:A�	� �%SRO:�<�_⳷�� �{T߈ч7x�#�z��+��������3�&��{u��,������c9�*
L����Au[k��h���G��Ŕ���s��zWW\�t�~�z�ƾ�&l��=Q�+:rr����8���/8�"��ڦՈW[� ೛�7���3J΅|��ώVd��vS����K�t&�u�? ����V~8<uu�u����Xs,W`���9���m`sظ$'�_o�Q"޾�Z<�N�/--ߨ�,g������R��C�x�p�X���f�[q
BD���x�4�ݴ,X�[�ݞ���0;s#�:�X߱A�}��v�^G�U���75����l�����A7Ј?I<&W��
���:����z��(� �c��x�S#Ϧ�Fl�j:�b�<ځ]��u0to�b>�f��!���zns5M|��v�*[���(ɝZ::�?�%׻����xxx�b��C�e�s@)	an�<���\�~��2�~8)���Na!Ҟ\��������h���}��^AE:���R3���4��8_A��萴vr�M�n4(�*��7�ȶkZ�p�$���)�|$r�m$m��%~AFR�Ï\8E�9�]7Y�U���:�џ{��v��
fY������wXXY��`�,U-ՊL���������]��m�\.��#-my���6)1	�Sگ8�l>_bI+ޟjܲ)�����|
�.u3n�ދ����5X=��~��qXFb-b�aʄ	B���mq���6�L��כ���*L�(tc���W�]"w/���?~�$󈧜vƁ�@{�[��6O=��ӻ�|2hSE%E�1�'��"��Ԝ��(��xS�~;����e���Q���x�l{�����Mxv���~D4��\�����_�k��-�S�@�h�i��D��� K�U|������s��Me�s;1���C�i_<yeI��r��>�q���)Jێț^ƻ�~=�N�/��6�}����3q=���[�=�`�!�.��*Ĳē�@'����P=u�s�EV9G��+((���pq�Hz���^�l����)�Y���$o<�]��5f��o�k�;�e�D�;j�S�Km1�m0���[rc��Q���2
�k;�C��^���~Lpg�0�dnn�,��8��H���44Zi��u��U��J����Q{`���Z�p�a�3�]I���`o�n*V�_�"ط�� и�����6Йz�oO �[���=��<�qOy��q�����S_Xh�Y£�H;����H_��j|��_��Ĝ���]YY	�s��A��omP<�!����#0�nQ�v��o���4������!-U�%�������:��}�b�_(7�U�C**h�Â�=���X݌�$����Nd9T%�گ�B"�h��rR�	X�O�ABUC��@'#���� �Kl�`]�v�h����PL�Bm���D����n���OT+�P�C({�����?�A9��upW9�H�2=�䈾G)���{��T�B�� �ł��>Y5n����濟����s��q��|�la�^��A f.���t��t:� ��2���������i�{]q�П(�?�;���ba*����90 �����a����hl���e����3��4�a5`3Ŷ�w�A�QJ��������'a����
`ʱ�+^����W�W=[�����g�

�b聹I��Bgh�C��y6����} ���qɋ'@���WXE������O3�h�F66�a��U�J��5��ܢ����ɒ���QD������L�L�߮;J�:dE�ue�v�5i���;���o�ޖ�b/��߮W�YJ(�=ϯY��tia�>dc�]^���׿w�ji�1�};Y;��VQ�+�^EB��x��D�I_U o��n0���;� {é�OP*R�`�l)Ը�Rc��T���-W:B�pk�ƀ���_@Zk��'�X���vVv��%�WW�Q�[Q��r���`v4ʨ�0ޭ�˔�t�B_�"n{�z��ث�.N�'f�kUc�����
N��֯K��aC���	������4%&&n���)Z�&��N��Ռ��ñ�X�����6��#�\�?���JI1�5�F'��������͍�ܒ����2�.D!�K����E�  �k�f;"�~H���'�kuO�jV�T��ҩ��1�q8?�֘^�ȁq�r����[����a����)�X��+�0�p���<�h �m��{�4�L x�'M^�	[���|��l.|�:�5J�ihb���`-�ӌ9MU��Ý��J ezU) ���|�={���]"��[�|�s7��Z�D��)ݼ�|:܃C;��y�^��^�̋
b�}�X�DY�mE{�sK+���.���=��y��hh�yуҏ�hc��H��ϧ���%���A�u�B��c�.N�m�&͊�	v$��h0דd�DQy�Yy�9��*?��V���?~h::����x�9Xwg۴��Y��Z֣�x,���me%�҉:��E���Warc���Z��9Tr	aOE������w&Ϻ[u���Uc�[�M�rP�r�	�>;�m�2��&�v�7?���$�#��`�_�$�-��V�k4v�X!&�Q�CI�kT����1�%V6���-�(`������ۆFG�Pj�f�	���]�b���âu��>m �{8t�/�3�?'��CŤ p��yг����s_(y�٨R��l��	!]�#�]|}j�����\�{��Xm', G�=�6|��н:��LEђ��EH�`Y<�B���R"Wr�\R���v�K��	@p6 i��3��(�ͽ�>v��0^�3g�,��ѣ �U��ʣ���kk��n�_�F��=~A?V�A�C����uG��p�AS8��;��<Q�f�<�<�P��Z�$~:�<N:-���O{b���zP�K������X���������y����	Rń�
�)�aQ���
�����޽{ ��i�x4��u#�|���g��@R��\���?��o?�^	�&��4�Z�-��ݕ&��q�p�<��Þ�_}��{��7uri�S�>n{����� ���6���D�1V֫�yZ��_� I��Y_� ��ge�Jd��Y�U���X��Į�����Z�X�_���l���?�"9�� �M�w�����O�PN`��'�������T���H��J8iW�P��ԉ�^��4��E������4x{No�	�)~�^�^���� %W7H9l�SbV�J�{?�|�I�Cj/E��{Ɓ"ST����h��D���zR~Iɰ��ڥ��%H��N� ��e|P����%�<��5J�á�&�*mb.q<0�KO��&X��׸�+�$y{{���ߓ�$I.�c��|����@]9���P�Z�Jc��%��K�}�c����>uD_9c���
�J�S~ު1���4�<8�E�v�嵦β ��S�2d�j�� e�d�d�yG�
ٱ�bX���W�g.�F'/j���g>�ty��-�E�~
�o7#����
 �AT�(�@x\��	�S~zz�{�_fS�pCE��Tzf�=h;$��OfųM1f_uѷ�v�7E����� @���xE:��Vx`ǚ����� u23/il�ߙ�
��X��#���Z~�4�4tt��i �GFX��4~2<����Y���Z���߅�^W;�6�.���v~�Gκ�-\SasM��Q�8W(�ĝq�KxC·'�Z��,��~-�gs��,.�\ۻ{hk��q�O�)H��%x�[9�(P�Lm��e����mݑ�T��j��ʄ<Kr��V�u�f*
]޸rV<g����M擛�98�ʣ���YO�٩�u� 1I�#��­TW̣cc�B?��\�*,޶��^nַs<��J�a��3��)d叽�����R՞I��S��㩥�{�2������ԣ�����!H�n����Qe v�OII�n{�`�ܨ`V�iG	�@)ł�M4�͓�������-s���tU����L�0>�ݱ�Εm��x))�����ڙH袠dwyq�k�r�й�[���L�@{u1���mu'I�229�lu���i��D��JY��}��#n�#�N�� 뢾�M;�HG5����E_����~�����Ai,|YJ+B}>�c{����[,|>/bf�O����$=�VP|"�zl��`cﻵu���3��}?�����_�ġ�b2�x���sth�E�\����8~v��$��GB��8T�!�5�e���E6��h����&cɃ��J�M�.�X#o�M��c��5�.V�q~��5��n���|0h��T�n��Lm\Ȝ��2z��F�gt	#����Y��1��8t�����o���k�/�`WV�&W�?>?m^5��� ��z�d���C`>Y3�9��*�W�id���9:�ߋ�����į�����6V�V�+e�M!9�5jt���X����9�?�Ф�����#�ư��7�(	�|��C��xmF�]�ӝ�.�JO71���lMF	2�����T<0nq��U��v�1c�ފ.W߃�����Om��o�Cᡫ֒\��5��VCe� zoYsss�|�+����-��䁻8��4�י�#I�t������z����|�����7���s�e ��Γ'㩱>^�y����C�^E�R���|��C��;�]�i��n�=&e#��HUGǊ�$�x/���㼹�9���e��PW�ω9�9>�ӚG����^����Ο���WĔ�?l����سtgɊ�F_��5�"��L�2��C�ۄ��;�d���Ӄj��Oҿ�bMP\̑�σ�����������v ���Lj�El���4�g� ]d
$d�F������2�K�1L��K�-_��� ����0�3�Nߵ�.�mZ��4�d�\�D>���u����$��xhZ�9�Yİ�+�>����{�NVtT�#I`�������#5���;�ѵ/��ĤY��W9�wV���j�-B1��CQ_��� o�=�s�_C�[�Lt)�Z�4��~����[(5����l� |�Pc:�q���V�apHǸ(�`#'v�9"NF	��u���`�R�N� �:g�E��ho%�����ŷ��z��b��So4�q��IJzM�K��ߦx'W�溱z�����w~��>�����'����d����y�(�~Iy�'��O�]�#5���D�%�{���%A���m~�İ�W{�\����l���A'�tC�0�Io�����0���Ϳ �#6�t
23[T��[Kcn(%����>D���r�p�"��+�2RZ���������!]����7ϟ��@E�q: /���)�?MN^a�q~i�b�R�eveR�kZ��p��8��n5�$O^$�u\V�F�:��d�J
������������뼵[��-���Zͬs�_����|��"G�D}rS����ޱQ�9u��G�����ӠZL���*��|�F��4T뉖��ؖF�����(�
������r�#v�с����LPm7?'�A�ؼ��K��l�>b.��b\���Z�,��� �Ed�v�E@��k�j�LK�fư|��+��E�B,m^��8,��»��j1
JU�;�zj�7�0?��lJ44�)�Y�p��>\V����s�?����u�9T�1�΅*�PlaY4�(T&t$�$��
�^��i�&T���S&RAס^t�^|lo	Uu�^��S�ӊz �!e=7g�R#y����p����7!-EI,��Xq$���Di�'�Y�L���6,7[4cטF w�bXf�å��ӏ�+d�u��;��䰸���'��U�<>����h�):+޵G ����E88�q�� �,��{�Ms�;)�����N��[�C�U9`�{{�Q<�dO�>�^���X�h�OG�VE�H�L�n(�"�,QEq\�z5⩊��~�uu}�V;��1ӹ��A@u���~�����V��}mʠ�zê�ZUk�ݍUjs���]
n�k�75�mU���vě����ĉi���9dco/ #c��AK`�́X�+(���7�q���lv\b�S������܊�A�kV(�@$9�O8m,�5��ݏ�$�����+�+�l/�'J͌���^?]���v�sc��Y�i]� $�)�ݸ	!s�P4�nx)[j�Do��.ه�>\����&P�v�I��K��*�Ҍ�e��e�B0hog��\����L�ih $T��\���y��VJ�q���\�Z,�@��G�x��㣳@��o�F��=06��W�Dr=u�n���6{�bbرf�,ZIac[j�2�������ht��3iQ����� #��W�6��5�u7{8�E����V�7t&�9�mʷ5ǿ�<Q�����]��iLܣ{u��ٳP]T[A!�o4H��� ��Ĳ�ƀ�;������j�t ��3~A[M-�P^f��S �5�>�w�}I�LN�=���P����fck�;�a��q^Hl���>�]���F�`f��|��F8��l���/J���]ۇ�֦�z(���۾�|G4}��BWn��S� ��J51U$f�^��ɇ�����5�|����Y���A
��e$��C�w.Ć\(�&p��L5�ڛ;y��}������,U�/�b93�Qt�8�<H��M.,�� 7����$��S�ZD�NY�O֮���lTgo���D8�$�&�p�ʦ��]?��<�D�#=��UI��`:������F �7��
��<
��x���[UME�Е��2�z���ϟ�⃙ 3��%D�U:
�O��!I��/fgg�k��Jj���������PI��ڏx�i�ڑc=�ު����d��v�B����,$����O����0+�۬,����7��v������{�I�Ц�P�|RX� c��V~���Y�*�3@v�;��2։�"���а�E�XS�	��NBe�Z\���G�E���S���e@�&n8	d�m����������xXa0]_��֖�p��^�K6�%��k��t�"y�N[wߏi���W�{����:j[�L�x�QH���<z#�?E�*�I4��`��q�ߠ�e���}������15��E�g���U�I��nwI�nC�Zӊ#v����{�ɡqzM�OV�;\G�@���*,��QjW���z������(��v)[`��ٵ���t�w �דz���;�M*rkR	ijB�c�Fc}�O�P��0��S��&D(�bf�߼gn��g��W7n��m!����j����D~c����%Q���@�R�|y�t��=ty��{�z4��0$� ����y��(㬹ߜ&���OC3�8��ǝ! WP�����T&q���"��_�� �.��ģ���]#�nH1��v���g����!�@�d	�Bz����$!G�ׯ����':��!qxR��:���)U??q�ۤ��Y~VJ^��bN�����ySq=Q��>�Q�e�2ν)����vpȜUWA�"��u����"�j��]8�;1�Yekn��{W��Z8h�i���! S��kvD�^P�+:�t��F�g$���H2 �:�Dݡ�%t��Ǹs�:�����n�m�GAqq/�Իh[Ԙ���P�C�	d?�K��H$J��PH�"�o�79��]�K�:N?hO�`�S�pPS�N?\�h�]}�^�Xz�����F�v�pO�5��+�l��Y�+��Ȟ��6d4߁]�G�hj�%�9D���][g�z�T����ד�,�̝���ͽ5,��,�ږ-c� _n��Elj>V���P����tu��/��s�HE���=��---
]���HZ��75���.0B�FFŀ�A����������}�~��2���|�}�*�q�)\���}�-��[	 ]K3h�{�����p���ܓ�/Y�+EzVTw����ј�h�T��z� f?M��C���o�.�ņu� !c
��c�GF�0�{w��
��L�L�
-��a~����
���3 ��!W��Ư&aU̙���!l�������M#1a�LF$+v��S�LnE7!!r��J|�V8�e93B/nG~:���P?6N+��U��%0�?�ajCF9��^���y���\�����[
7�O�D$��ȭt������@�҅��C����ᢪ	��F4�_	�9&;++YNNN�i���F	 ����e�� �n�8a1_!af�Rq>�S�R�<���Lx�f��0�5�b���e���B��7�2xɭ��Bwe*�_fMϮ#�U���ʟ�&(��e0��9>9kJՠ.�YE�x.''��ߥ׏�C�uE��SP��Y2jt�~�S(6U7�J��������THv�R��S|��4P/^�nN�Ra.���%��Y�������ʟϋ������֟���88����7�{/ 9�h�m����k�m�o��+�r`����re��5�S����c&?�������Z-����%�=����ȼ>�����/��^���zhh�Âo?b���}��I9u�˃�~��;. �?�'����A}%�b�xJ��+��#ԡ9�I��ݴ)go��d����'��<��P�㥦Y� ~�Dv�{A�G#����Vڵ��y��ݷ]}%_~����l�GpzbK����x�1`�.݅�K� ������֏�L�1h�<�Z���#�x�r�;���l7�WN�.Yz{_9��m�%�2��Pű�[6{}�#*/S��2A�r��X��w�^�-������ȉĿ�:Y	�e	����i��^K�~�۷�l��U���$����:oa�f�
m���R��qR�Ƞf �ݥ���0��|�ug'���'�Β]w�^��.���0����Ǎ� � %C�b�<�{�8m��w)�@�`Re�L������Tg�l�E��&��#�Щ/U�&<`�X#̾5لڅ>�z�j�4Yd�2�N�|6���crXhߺˣ`%��d&'t����.A��5$޷mq��"�/t�!sv��]���i�JWI/5{A��-�⫛�� �۴������������5��0	h��20;�cş�%���k����P�+��h��v7]o~ɍl�c�a��	ǀ4?���5����4��� /�b�6�7���lP����nM`��p;X
o�x�7ܕ����f�����K�n;,l�m<(7؝}7�)YuDZ���ɽ4��e���RdZr��(b[G�8�̈��OE�O�����t%�5��#���c�H@PP�����\;�v�T���ں]��}FX�
��������z>��.A�q^(�y��.�&���7#Y+2���}���Y_�c��r�Jtg��_�\��ߠlo�Mv�����Q�G����/���?mFI�Q�8��=�FH8𝛇GR�����B�|�S���q���á����}l�c����Vb��B�^�\������̭x<�`��g��͑�Ӛ7�A��Hp�!BI3~,E�ѻ*������� ��@�m��=}\�����H�- �'S`���� k��S�^X�.1,����;]����MT��=:�*�=���5�E��.7Ut���.r�XS'�ݍWS��i�E��d����u�T��-��0����{��h�݄-��&�tgi�O�T�ƣOa�P�/{�N<�M��A]���-*�A��	LM�����j0B��
x,�Αdu�zQ��*z��γ�׻q��o��
o,�{k~0�ڸ"�~�w�+�jdz�j40��/:��*}�V?�֞���D���Ȥڽ=r�GrK+�m��91v�G10��������I 7�/?��l{y S
���:hqU'����'є,#^���c�̩g�_�����*^�.*�4��7K�NDA����l�$�k�lq��E@�=�H�(_� g����t����c����h <��4 sZO1z@�	a��EEE��W�**+���Q=��80,�������)�R����n�����,k��T���>-�	%[��G2���Y8����r��<7H��b���5�U��)�k���i���OyHmF��+@Dˮyݜ�Y�����uh��R#��Znnlć=�[�04��wV�����t:Di�[���������<K�?�w>�9��9����5>�A��c�̳����G�Np���p&o�c��_��]�p���	h�wT��\�ؿ&>�ŅQ�_�#@=��KwPEf��r���X�!Y�UQF8�%��=���9����ٶ����N6�=���W_��*�?�	%$�YRD��Ai�X�DB�S�A�C���i��]����"~��^?�����Μ9�yΜy�Wgp���s�Z�}G=��NMv��)��K�J��8J\gt����w/)�o@��g�q��cD�7�&����}e�2�`��W�VHF����Y���k_�?/ѫ�c"V��6������Oę�PR�����,'x��t8e�Q׻��G0�ȫ=d�s�bmOً`JO=0��y�V��oB��=,)�E)Hq�z�IҫH.��d�m�,��hfkcm�}�5��~5!+�����9R���WT� ^��φ���P�����&���	55d�R��tX� E<�|M�����
�w��Ԟ�|z�Ĭ���'"����$�}��뎞�#W�yπ?2��k��������'�ɷ����l]�'Ǆ>S��.�;U$��帉"Sv��VG�|��2�vh�w��ߦ�8��L��w��~�Gt���TW��)����u��++G\Ü��	�@�Q�*�U���;�,=���ja+X�Q�(�(��H�ȹ'�b<����1��'�������D���?�-�T�x9�k'��҄���}i�~Af/C��׶��n�6���Ю�F�y�d��㦔Wb���QW-G�Hs�g�i����<:�Dz���Hs�b���M�Ν��;F���
%2WM��Kݦ T\s�4�$��JZ�~O�Ù��k��5T�ʁ�©�DL�`Cd:W�cc�z�4�2m�t�i˄`/ ��tu��q@g�����<�H�U~����l�x����\5 ��M=#�Nv��,�*`ד���/3)��:zId�z/��i��~}�w,������6%�'����w�1���is��$�uz��.�/P<�ƱLw~��(;;�	�:�v����<�0J�*y|k�\5q��҂l���ד�21�`�K33�mJ�Q��i,%��O�k�-�&��Qrp��ay1$�;���u�/
�gy�M?͇DҦMq����{�!]���[r�3�<��$-\r�*�����pnJ[�`D�Щǥ~����x���{��̓�������h����GR��kv-8�@n�2)�4��uϰO���T��Ȉk�|�S ��'2��O��XܾE!Y;^Kn$����I��f������PWq��M�(萬�� ��ëÊL�����]o��׵rx�l�kc���Hx��m/M^~��M"��w��"����h�Mk���g��N�3�^�Kx�*fR�q�YX�Y�gΝ$틝+{v�~6����� �sC��cWAbx �	tQ��V�p'N�W���ٛ��P4��+l?�(6���n�z�6'5 ��^�]��i-�6�g6�უ��j.8^���\*#>��Ǟ��2�Nֺ�g�m#V����\���ù'���=~��^bXR���a��3_/,(�q�E���'dfV(�ߣH����b7���0�rƈTy{H��B�C�Q.ͼ.P��Sذ�����i��<kn��� VOU�5kt}�U�"J��z�`�\C��а6���eۇ��#���Z��y��,`�-�ef��w1��y����7D�r��o�mt6� Lr���<�s}{�?�3��A���]�i'�fӲ-J"ojWW���҂Z��;��� �`���NJ{k����d�?���Q�XIOBJ��ɞ�K�6(���b��n����[�#,���:�--6�5q�2@�f�jD(��tMhyu���M���� �d�}���*o<�
Xcf�E�L�B��,��������}���#��O>�C
�v:|�g۷�E�� J"\꿧Ֆq��ui�kx�J���5?e��p�;���Qr���-�	���k���+���^Ű��g�F�V�ԧ���)��(9���$`���؆J�L��s�ز'�H568iz�5�{)��̺{������8�����á	���)O�QY�9��6ؕ�`�4[y8�ΒDy3�o%�.��.ץo�b]�^V8��3�:���X�x��V��=�_�|T��xg�WflSě�=�xRte�,��c�o^~�Ggr���X�UJ��}i�;�R��� �N��E"���&h�T�%˩�-�8t���d~�/�`P�r�'%�M,���S��-����B�d��=���az�7������K��]Ǝ�8�f�vP�%.�;$��֜��?W���k���u&˩;扟m�b�&��Z�|^���aeeb��M���4���5�k�`v7R�7<�0._�de����2Q��8
��e�ŭ�6�V	] ��n���B�3*ؾ@{��n(8vcT�B}=�ۯ�x�����˂C��v�5nypK��#l����R�\^yGB��mʻ��^�o�#�؜W�}��掆:Лݕ��Z���[����(4�O��F8�Ngtj�8B�bn��2��Z�xM@���� ��3�t�,H%'^{���駗������mm�S���4�ͪ��F_�?wl�j����ޑ5c�0��O�7g�_��u�<�]7Z��;��bз�b������VC�O�����.�������0Ei�5}���t��w7���|�qά*����ő���+�<�~A<e=l5Z��^����K���^��g�r��b�9�M��g�
����}pbPߟ�?%j�Os<�
�(��L�di��E���3��؏�Bஓ��l�T�,F}2a���!�_���/�ȫ�R]ΒC���N6%a��G�����I
���w�XHC��� *;"�:;�i>����+6�ʻq�:`�9]Դ�=4އM���j������'sU-!]ָ�f���K��5���Qؽ���@������!0�C5f�m��ڦ�Z�C��SS��o�ѝ�(�����+�Hkf����	��)���x��^�6���nd&}/�������I��I���pv��V`r?�aJT�0�����W{;�-�;�c��
���q��'��<�rO�e�rUMH�'kr�T���^�%����Ǐ��Q��A�.�?�Q���Յ���gs��ܕ6
��H�KP�c�:n͜X�͉����x�����Z�f���Lja����9�����o����sF����=خ��Jy�e׹<?,������ő�A�1F��џ�����~[ݦ0��C�D ��6Lc��#��X����j1r� !1�Wo@邏����ݚ�y]��/Vŕ[9v���dӥͨK�ww	�����U~�I1�P����j��7�Q�x�S:�̐�7�r!����'ۤ����n�ov��	��*&7�T�d��2#����{�Ħ���nX2��0CI�R}0ť�k�O+�Z��,L����V�%�;�R��-���SL3эv&���R�V��J���(��:�w<��E킻m,�y��-���Z��C�7'��s��p㏵���>Ϣ�9X��d	�0�)��&�
M񮷱�ǒ�I@ۑX�KXԌ`BeJ�����.^�Ձ.rO���L��,�}%k3vύ��+��Ϧ7�w��OT��P4�I�.5������>4�2��Sڤ��[l�:<K����uK�kc�Y;n�u{R\���md݅Gs1sb�d,�6l	��:��U�{��
5�תTT!�'���,�m���B����5��-�C!u�/��=���4�����mK�_�<.�*M���f��.`�iƱ��K-#*����y��3LN����~���9&n�X�9J������O5���E��4>��By6\��N �r���SѢLq_��]cl`w��Vz##{�����	'�=�a��;���]{���#V�TA�,�W���1���L^	E�K'���0��`:��.�:P�ۧ�P�~,s���\�b�~�w:o����-���q��w0�^H���s�^~��:jb�^�?
�h���V��0c�lBccF���g����柜S�w���&l��z�(��g]���8�T��i=5�O���V��zs�?�t6/��Ll��<�'3����A8�<j�k<�d�ږV��u�l�.�4tV�(Z'̎I�_��>�8������,��K��vv.8!nu-970��eom��e� \L�$nP*r��(�`9i��i�q|y���N�����Z��u���'/	r �;jT4�R���i�K��G Ŧ��o�R,�Y���
�G��"�nb����N��o�̓�i�,+����>�Y2�Y�6	�)�u'X��@	w�� trp(^
aX��c������u�Z~�L��ҭ�t@������;�n�yiDl��l��6
���}� Bu��(ؾfS�c2�~E@������:�#��kyq�`qK-l�_P���������3��<r���Y::�~�o�p�kQ?
�<�S��<����W��wF���|�B�7[�:���1���!��#[�0|-�\�kv$EL˥99�&
���CT�j4�)B��+���7��^u���#C�3���6Y���R�e.ڟ�l���d��>�ĺ� 
����Y�(`����J��ݞH������:�Ɇ>�D�2w"�VEf��R��ѫWG�'�8&?�B�.=>v:���ȑ�i��ƻ�Z�S����v��m�c4����N��{�<S����N��y*?�9�G86�`ѻ �B ^Ƿ�@5Ns�5~h��V���=	�*|�O�Ǔ�w�(�z|@�Ǜ�rP��[{e�88�B	��s�0
�{���Z8Q�Q��$V7U�N,0.(��}�v'_���d�ϲ-g������kj�-��g��������}�.�V�\����bN.s%�Ae��)�F:���%�m5fkKo�'Hu�{�~1zZOU;vL�A��Y��p�|�P��fs%����Ǽ�|x�נ�Noo���Wh�������S�8�j�|��00�	xy
�'*�g��Iw����	���@�����ox��uQ�1�ۇRL���cP�����zܳē�5ν*@���� �.v+'2�/����.�)*�vh����Ǿ�j��d������_�ƫ	$��p�e�V���.�a��rP>�T4�ш*����!"���|��F}ҝ�Zş�������^��RXq}��R�zE"<�Ok�/��f=��⮗�������#��X�M㧺zn̜�h�U��c3kȠ�*R��x��Pt�$N�����/ⶌ��]�ё�[�I69T�nc_�p͉y��	Ji�ȋ��_�0�>W4�ւ�u.@G�`��4�3�E�r�3Q�T-v��'�%�g`��ݮaN���6����+�#�c]Z�Z!9�&��@X�bHhi��$K��}{E��U�B����6)���.��>����n^�s����k�����R�D�c�7��&j���D
N�����^VC�:�
�F��O��^�8�X��]%�0�I��n����w�ݓ�p�Q����
*�b�4�[���Ӝ��YSD�'��+Z��kQ��*��R�y�" �����
"Ï�{&�W��湄��V�.�@����	R"TK�zb���QP����7�� �^��j�G���Z�LG��Qou~����߉h�">�I���C��/�w��*������� $tO�]�P��^��<%��� egHć�É���}c��<�(:��#�R�}D(���HA���ø�_�~���3P귦�XR��g�{��Y����������-�*C�w��"	K���T�ˉ�� �>!��N\���f��3��s~.�-~�(a}�"��ܚ��^B���<��		���)��r�����~��Þ�~ s�� 8j�	Q���;v�6��"���y�zOzWl�-���&��]��>��1D�[$6�܌JR�<`+s��<[)�W�G�\C4����;ܫxe*{��fl���%H��;|���A4~&���,li�qC��ظ�n���tje2vf樾8�a������ɡ?F��|W�kȓ���h��6�ũ;&�	�H���~���Vj��k}=z�y��/ʷ�2}�J�'t��	Ҟ{ T�0����>0��M��|�G�~�~�mP�-k���g+C��BƫR�ǧmyy]�o�{��m�Qeh�z��Oa���V��jxP����r�Z;������ܕ���OEo�uqWS@�3�A{�H����8sFs)Om$�/��aT�;/o�������c�#����JL��c����P	��ZsqeI����Ζ�Aa����b�w���(��=�D1!أd
ʇ&�-��/r�k+�[<��G��TM�n��zG�Z#p��+A�6n-ѫ%������Ye����<C��T)���w��E{�� ɓ��� �Iu���É�XV����J��l�٬���Kq���/��E���]	t�('c��7�kbYY5@Լ|劢�`���܎���î����Ù��iaiJiB��Qv><���wG�Lc@�0s�t�%Aۃ� ���/���Er]"u˘��]��}�S��U��V:y��g�w
-'�ߗ�R`l�om�ޡ��8���F���Rt����)L}�+HLCU5
��ad4��J
���?d3tLș���#�f(���k�N���أ���>W�12\١���3��O�g���qU��<�]7t�\�H_�J���U���z���t����G߇=x w#��H�6O���+L���m=<���o߳rU�>R^~����nM�u3n)h4ZA��5�9�*���&�m��]�腕'���h�Ј��C^aᒑ5������li��;	�6�;�9Ɖd`����)�s5oY��q׮�}PN�M�z*�!�E�Of9����N�:
+�����L�-����=� 8Ȅjk.K- ����r�󊒲������h�-G���6KY��O�~�U~iV�C�?�B�Gg�[K��W����S��,J|��ɑ��i��\�o�B��{'=nyyy�LSUُNp��3!L��/fc���a��n�Xm��ɋ0V)�8.�XX�s�)�^W�tI�q��ɸ]}43K���G��aBhhF�n������b��R�wC���c?��񂢢e�-"�]X���|�Qt3��8��F�n��{�<s���f�s>�l'H��>f���ي���Qܽ�M�vV�rg<�I$�֝HZ��p������b��a,qrޤ�x{�o\7��ɍ�8�ʠ�zX��V����@���g��_ۻkB+LC�}��|��� s�Y�5[����lvCL��R�wY�����o��������$v %I��ξ��.G?:\h=rFID#Z��	����5���h�"ǎ�f�:(|��w�����Lpf���-}ym����\��`I	ｵGT�z���[ʗEm����pd��[��[�X�c���ǿ�w��������5��&�^�NY�SR�n\:���>%W����^t�w�(+5}��13#�(tFݪe�;��u��p���sؔH��KqCXņլPW�"��.EÏ�����?�%Ɩ}�l�����*�R�Oxdf��'��"��>K,���|<�.�|Lom=�
�
q�>���{(��7>���Ւ�m�(@9�v�Ѷ�.\�O2�u�/}���p*��垞�V�N���Y����/�O��ygy�z\3^�f\�_�G�O4e\�t�n�3�j8h��C#M���;�̥D�NR�A�6���YJ<^���|�	gTE|vS,�E��.��$���m3���~e��W��/m%���c~�VlCH'�� ���6�t����Bŗ�$aVy�阯9|�%P8�������B��1Y^����rD�T��FN�
�����.�ܷ���1�mz��I'>&��<�5�t�\��`�ݗܬWՓm+�f��+Ԛ!4�7�W��s�챠5��o� 4��]�`���-~�n\�ck��dm��Jt�j0��HEl��a���0gݶA��_Wf�0������u�������X��b�2:^�~~��h#�^�x1D��L�&�����C�PX���b3j���A�ռ��Pw�aig�z!L�06�Z��r�5i���)2sJT�����ntF�����C��ABy��bܖI�<_���<�zM߳C�c��E8b��i�:$�!y�Dv��[���+�6ϖ��t��ᦄ���Y��'XE�aS��o�M���f��� Cfk�w�K���jb���WQ����X���܉pqM�_���y�@Xm��
���H��{�$��x�N`lF,S�z�=���/lmG�S�>_H�TU�_>n��z���I~Dp%�.a6GKm��5��m��HɆ_���K�o��P��>11"r�e�s%"9I��t�i������&�ΰ%�a&-͖�%k�m�ǎ������Y��/ x=��႘�='a���Ld���\���EȺ7"P����"���?�=��=��-:�Kg�^��6���9^���m2F�o��P8��\�+';XtI�Û��^��:�Yg��%���M�j�m�g���8�I	6���9X���s�2N��o�B�Q�����ņ���m*���覾�HHI��et��ɍHs��>�suB����vRc3�n�;f_�#��͔\«�jkD�ˊ�������V<E�06�.�$B:)��F}~�3�4E����P�b�;#cc�K8�h�tS�@Y�(����-�,7���jg�t����N"�9I�׷�7���z��b�S5\�ss�a��ϼim�q��bB�K��\n���.�fU��O�U��s4q�bk�,}�� .֞P���L�˯[�:�e�8�m���Vz�ڣ=�F���qA�?h���7~���iC��W��O�B5����R�*���S����`��NNN��ЛU���x�f��l�� ߤ%�	zH��z�ߧy��p���M�j!֢?1sm�L��'*q�{EO��f)n��x��S9?��C�S��3�z��Fw0oZz��.�(�W��i	x��s��=k��i��basG��q "M9��Tۄ�%'S��U,�ޅmz@����k���cd+++!������r��pg��U�T8�_��B"�p�'�q�O���iٛ���`kr���$�I�0�	>{5���yG����nN\��/�3O�k��}@��D[��\=��V��S�G)Vr�Y�����C��'�[� �O�J�Btnmo�<�]�V��N$jiO�>�w�S1�3�q�Z��Ҵ��quY�:�K�zl�����{sAK��˼#7��9s23O�9h�F��ϵ��ׂѢ�P���7ta�7q�o3�N�3������{��ш�΋����FX੣k��)����M�ou��E�S/�F)��A"K�
-Ặ|)��IC�`|j��,���Bֵ�A�W��d�b-�W� AĖ_�M��>s.��RF�`9�Z��,L���ԯ�h��z�r�=Tkn7�:�fz+�6X��������4�'z��8�A�y����R�������ZҟN''�� �*<$��#rn��*����Z���(�<�H�l�iC�9�J����Ӹ���u������3�13�4>=�y�q��5)�^��Ɋ?X�!��0HV�>����/��gff�R|��K�M&�ʃ��\]G�L)ޣ�i�=,	�=�2=��J���0!��p\�W^؞�V��Gv"0[8q��`^@��L-�#���.�@�_��'�����\e�2]H�a�O����h���4���]��څdK�:�T^��ƍ�vḷCB�/2�E�-��i���y�ڛ;-*��p1{����455��J���>j���`��~�*$����Q��P����K8cw�JY#[0B�K���o�fjj��y�<��P-^�1���f��$'��^&ك�!��V�G���8�GGW����o���� %��-9��oO�a�"�8��|��+��~�
?��@2ZV����b����]��Ǜ�K+]_�XX�>����L�އ��^�*]��Hf�����GvrQ2���T1�$dd}�u~����/�s�=��Z@Vp�%.#��l��T��=8����FIB�p�{��f*T;�Y�r{�F���ж֔c7i�2��[�̈́R.&�i)Vƚ^�~~0.�\P��|��?o����"�ǧOuс�z�2	|[>tpS����:���0/O��y+$k8�*�˷o���-�$t�s{���A�7�B�[�=ys ���r;��p�����]t�l���D���AK�ї�M�hƪ�܀6JEZ:(9%z[�?����n�Zؚb���D>��塳y �ڮŦ8!��p���\���I+P��h[���>�8�`3�q�W�aդ$��͖�	}ʜ����=����o�)4����_��g����\ޝv�^ꍃ����F�i��+���I�^��C}��
�l�xxV�+^���|Ms$Nf��;t�0�Y��=ٞZ���;/8/�q�4��s��B��Ѕ�<��&��G���џmMCC�񵍍��b��,���Sر"������nk�3}�t�.zh��4(N;������]\�=�$���ƥ��M���6ڊ��\�j��{Ez��nk��KC�������<���x:�q�}G 0:�v�Q�$�j�B���� )��=7D���Y���rr̦˚,��h�:<^pP؄��v`6V�#�y)�r}�w�h�M��M�I $EI~���X�,��<t UP"װ4f1VRu��pJA�u�wy�V2�a�����}x�@�
�C�x�Q4�#�lS>�_�y�M���Y^�m2ҧg��$���=e���Ҁ�i������>�H$�-1�G�g�x�"��d2�\yۓX7�FgA�S�hFS[;?�۲��^��Tyv������������������Ʉmmlz����f_����[���+��a'k��w�@�E��=}�i��s5P��6L�8:2µL���B�cR]+`Rj��5�����D|�m��|ĹYF,%�`/�n���.N����j����#~�Ït����j����Q��P���2  @�.�����5����bv
	郍�;4�������¦t"}���|�0xX�8;'���Tk�>*�?�9^�˚���Wv!�,^���r�O^\)�·�pB����R���xyye�5TT>|������`x�T,�A[|��"~���+�:88 �&R��HPP��q��w+ ��PȯN�\�r�x�W�{������˭**-龫/8�wl��0�T���Nc������{��> �斖�YY�G(Mwwʘù�֬�����+<|��m^��	0?5� z 4(((F��0��2� ZW(!��AZݲI/_��  С�p����T�|�j4ONm-X��Җg�>�	~���Rmk�4�*k��b�W:E3<��1�l������<����o�Ù����˵��F:��@���������u0�ɤG�oO��N�'&&�E6�#D�R�������|"[��'�hьA�S�R�t�V�*�	.���謯ܤ^4���N[���؞iG���a�~(ƅ��s�n�����)Վ�낪��u��	������W���V���!�[>��L�������ܐ|��+!��ɩ)H�D��l�ܬ,�P2�1�wJ�_'��`1�j�	�x]n���N��&9�q���f.bv+�+���J{���5μ���S*��0�ȅ3��ӻƣ[5{o�9"9'8���WwY���B�%H�LSCC���<��3�+4>��Lօ �������1wr�A�:�Y��pk���?E��M��f�=����1HU�d9y�����n�S�߿�=�&f�U 8~YP�Ch#����H
}F�}�x�2֔��	D�6���|"�{)��o�����o�
���<���F0�еsx�5�3�w�xl���n!t��1�萸��CoŇ���څ���K|^5�
l��AQvvZ�N������'<gJ-iY=��;� ��yKO#���[�Y8���RfK����'þ���%]�w�mf��o�y����쑑�3'8�H��^���g7|�͙���4��(5�Q#�^���yy�G�:��d:��{�	�*E0�6��{�K0v�#sw�_�w��;/�d�z��`"��Ar�V�h$3m~�
SN��a�xG�-��uHIz�'s݂��2zO��^Hɇe6� ��3�c�{H8{~�Y�B��|D! �*gP�<F�5��{_j���8�@����"P2A6�bֹ�,��5�b�|iVś��[pB��Qr�'�27���7*��uT4{O
�D�x���ɕ��6�'�c��� ���g��qr��C+�(OH��mʎY���&4���%M>����d��j�WiE���K
�.S�7��PL���8��ۇ��[�gZ��n��1�����·wh��:��������L�P��o�3��� �ܫ����;�b�;�Mי���n����O3�������&��N�y�)���}��^l:Q�W��$Z+/D� ���ޤ 9�ΪO���}xi��ۺߢ�������h�x�}�RF�/��9>�[��?�4��C=�S�p���4�-��܆pX���n��/���DŦ�:Ăg���� zB�����TXJBHq�_@V�*Z��[Zyj�3E��vDw�Ŧ��G �z�r{j`�g��-��%�-���\W�w&���Ҁ�8���Cwg�#B�3�Y~�)�r��|f?�����O˴)�������{� ��P�T�Ҕ�m�ȡbO�X�z/R�b��c��{ͤ?�Z�h4����>���}}U`4�6W��j`�TU��;9>,=��� G/n��T���`�`�]Q�Ң�3�Z��4s����������������!����|�~�Ը�˂���{ISM-z�e����q{PH��ȌR�`����g����PN0�L(�~jo_1-��u�ζ��;~GC��#!Ε;7iJG2J��ˑN&�Saa�3�]�c�w������82��BK����Oթ����9���h��p���.�l[7�>���x�ծ��55Hq���+ �iH�5 yBK^�up���g���FZZ�P�"Y��E�'l5�j%a��c�����fݿ��Pڎ��"}'1$֢ݺE������72�����n�ś9�>�>�i8��B���
�e�"@	�hޮ�c�vT�k*���u��,߇�f��L�$�1�s�!�����=j�[�L^�7V�Q�J ����É|�Sk���g�����6:��(ࣷ�{�����g|�����\ /���K;��AK�zz�9#,�& ��.g��Чb^�$,թ�%e��I'�.��ׯq�0� )���s�K	dx]�U��폊)�D���R�;��h��^^��~��HG�F������V�X$ �ɏBUD7�A	F��R�	>@�x6}�����z���m�N\
|�ZWp"ɡ���I��E3)rH���W��g|����!� 9?�6������cc�%i��Hȳ���X��>�ՅG��]�����\Qy�z$W�Sr���#b�Y��V�L}��B����U�=$N�/K#�(I�n�mC����>$���k����Sy����ݫ
����--/�]2Ժ;� uK�������@|��zRq9MM5LJ�v�I�{oM��C�ZQY��VId��rv3�� �U�.G����qn����,n���C1���抉$���W�N�:hoA*��47OC7ůj֭�5�E�����'_�ЕRv��)�#X���-W��p�꺦l��[
��/%�`�ia#ԣQ{����Wu�e��J�p��MRR��!��'��V7m��CR3�G\����@X���[�>���O���SW`U��t�<�xX���tX�+,���MHD96�GŰ�[�� Ń'�L�����J�nd�D�ýX�H/\�
�~+�~[]�s�[���j�B~F�OD�逸��؊�ȓ?�lY�ᲃq成�=Qmy�/s�����55N:)w�B��yvW͌��z�vc�4Q�H��#iI'��5A�Z�W�6��{��L�.��U@�+'�ٛ���k�Fw��+�T�(@	b���9#T��f�/M�j{��*Z���������,=��ګI��P=���H�*���Z���f˓��^��_t�F��с�d��?�k~�h�<)ɋ�ia9,y�%S֮������n�m���u>��zӆ��R8Ru���1��3�)&d�~���Ց�[y���6�����{.3�je�V�}�|��@ ���k�B�5�r_��ӧ�HU���谸�S�7ɒ*����A��|M���k_:%"%�A~��6���ǈ��V��~[��N�&��Z��KIY.ˋ�k�'��Y�o���wp�@��ېB��x�8[_��q� �S���2���.�4����2w�p�f1��E�?KȪ��\ֲ�WS]��J��)WO�^oH��W����o'��V×��h�x ��lû�-{�{��}^��5�$�6�V����-|��q�(C�#gs"e����o�ΕΫ���s>���Eތ����%��d�G8<sg1����ߺs��b��e;C�����g�m~�j��ϬpR���4��<Djb�l�)6.n�~') ���]�-�G�����9�#XU�ü� �� %�����*��Z�\P�
���%�r�K����z@�v.h�`YYb�5�W�:sM���8[uL���"�#��B�V��}�!"�����?��������N���NM��a�Z�c�bM��]/��STbr�g-�2Q�:�{_m[��s+�s���+�4n"-uDq~�4�E�7��Tv�[[�ɼ�|)����1S�u�V�B�74��N�h���v���Y|`���q�u��[��"��᪓)��	S��0�{?��m��r��T#Z:�]��z�V%�����%^��}:�^��l�g�[ib\�D�֞Z���3���U!��.	6m�����Yݔ����ann^x��r�*����$��%���J�C�q,�E��FJ���BVn�S!�u��M(�FN8��o��[��9��؞H�#��O�w��Kr��٠�(���������R���((\	� ;5�R��3f!�JW^�ܸ�-�wj��-�g0+Gj�٪��ܠ<��`L�=�����A�D�%R3Ud��贺��)����@�3&�;��_��]>[�\?q�r�~�~�":Q��&J��A����t��=�q���jW){�zM�]���#:{��ʩ�!C�"��",�L%�w{{�f�k����l;@��F�����S9zH�h�uCBBx\�@\赨�����E[��\�9�[4�<x� ��{C�t!C����}��P;M�'֭�  3x���?;CtPf�ȟǓ^�(��7�w��W�|���w��t%�c��Q0��U��Ǵn���+�@�ͭ�/��;��}h�c&��v>��s!���4��M�s��	G)�e���iJ���ŵ�Z���1[C��F�K$g���.�1k�wx4��:h�`�=�m��ϳ���������U*c5��E8�4�w0�~�Q�L�a¸����� ?�b�t��a��j )��H��y3����
�-OʭƵ�,�EY�rɗ�
w�Z��5J�O�I�]�W4(m��ߺ=k��d8Fj�f����-*(Pn_�D'3=� K���4�I���u�\�����ESO���:@J�g�A�����:r�r��S��j�\�� 1�#�]Si�}���rߏӿe��K�y�t~����omu��^o���/��j��pPm�H��g����J�82�ͫ(̜�۫	[��)?5�l����%�Yk%g��j����ݴ|��{p";�O����f��8[gТ�0'G�]mE����qtf�t}�8����J��xxx��Uuu� �_��������ԧj��zL�|/2���}���>�&x5��sZ�W�B�g�}����O�EY=t�J6#���s�n���V�|�CF!�����Hq���.@*n�c�*��	ZliY7Y{�_H��|�x�ޔ�ib�eV��bI��N��M93#�4� �� _�1����mw�ɇ��._��#,|����m5!P�㘸�u�񜝝c�A�\Z\챐���K�11�tn�_�@��Q�!Y?o�����N�z����bS��6�[�ko��+��+���k�����Ma|�������R��O=�"��v��b��t�;�.,򮟚}�/1O��i�~zg$(���
Y�pG;XR�=����zT�}��Znn{SJ�=��q=PM9��!��'���	S�x�5c_�p�B|ݺ��
*���v=&������H�"yϨ��Fad!buX�{wb[��������@����?_0l��*����/Ūԉ9�?�ȋ�����H����o���Y*�*ٹ#���d��K��W�eo%t�{��$f�\���>��&+'l�<����ˬ�f`���q��/zc��G�cr��( �ⳟ.��Yg�-�&�ȩ��x5+Ñ����_i��)0���̾T'��%��'�[F���\�|��R�j�M���9��kcE����:����8�W/�����#�F��f�llj*=�Go.go��u#�q��qO=Pj��˻m~��r99��&�&�9=M���% "��vkE+N;o�|�=�ƴ��ѷ~s�uI���8�Ie��v. ���D�d��)�d��P������$�l��R���T��|�=��:���Z�^X�%���������{ID� W�����D���z����:����;Ϥ�v��zՊ�
�������n�Ր���������_pI��i����w(R0p+=]g����xJ��ԟ9�(�;g����Od#���{��d��W�H��t�=���"> �tʲ�_G=��r[myQ�]��[�����I��b>��N?q)~?������W�!��&���i}���7��p�w
cd�ǔ.U9���*X�B1�,�r�(�/{{PH�M���$m��*>d	�Pa�i���EU*�դԫI�S��:LW�,1����pÊY�0ӂ�o�o�D�6��>�S�@�GSsq�r��O� �͍'��H��W�͠^e��}&1�fP��ROdr�.�?��3�Ҁ:��Qq^�z��\q�S��r3o���25�c�wT�M$s����-�I�����M��v1��l��]�fKL.�֬K�e��O�A�d�����8�w` :������p�y4�������[��]�e�oO6�Y�҃fo�|�+��~�����/�2�r�(5TF[_|P��h��oб���� ��Qx�H1߃��N�>kk�DD�z/{7��Z[�K�+�m����� ��ׇ�6��"��p��
}ZyY��
)[�B�`�;���9�~���d���2��D8_�<Q=�bX��O�0��X�9��o?q} � z��!&�L��O�	U.@	�g��z�p	��,˙D���|7�n�'@��oD��x�x�ߝ�ŉ�ɯ�g�m��|�q�����g�����{;���U����8�jF	�"���1��U
�V���:Y'�pg�'�D�~U���=m~��}]�SȧUp��n�V�����¬��������۷H���]$�e�ꫝq���"L�=J��Jt�D��oD� �UL�{���h ܇�6��R�MW�5���o��y�*I;Y�Ք������N;���������mJp9>����`����<�
��3�v!�0n�n�1/��'��n�?̽wTT˶=�r�k��((�@R$K��Ar��AA���dԣ�( 9#H�"9�"Z�d����n~U��w����c����Uk�5�\k�]���x�A��F0?���B?��p�>%!���l�TE׈�l�^��w��*�!v��/�6��@q�x��}]xw-��Z��wD�X��^�#�$��CO]ͮx�H|⹚�_�_�N��G\�9K=�2�Cɦ�;s/�6��ͅ/�T��:�,ѷ�@K8&:w��yI�K�G��Sƣe	LS33e�F@(e����Xo�D��aUS�/����y�Ƈ��>ݍ�vA��?ٳ83??�� �Bl��+m�'��(v>�cYI'�>넫��:���������o` n���m�[/�T��v�\��:����Ļ}�W��d?��J!+����,Z�ru���͒��tW��N0D<̱,���M����������u2?�jxs��*������/��l3��O�b�e��(P��� J�jLM`��S%f�����:�P�^����ss+��iQ�� )�]���}2>z��9
6#y6�d����+��rkuOx���.6�\,ML����%#|�������
�����率cF�l�f���5��?��?�@���L�@.�X�@�y�ϕ�E��X�R����N�����Em��H�2ӹ�Wh�����E�N�P�����q������.{Q��1����̹'@��DK�����+��P�%���;]9���m��h����8�m��ҋ���n�i)-u�Y ��#t�G�<��e�)_֋�ݹψ��_����U���o��>��i^�ւ�m\��[���y�"�r�bq9�gMS���6�e_���kfq�,�ZMEW7��������)P6�e�����,�)SC��%�Ǔ�M��V*��P�;e7�[���!wsn:������ Ǘs�"g�/F�pk�GN����Ѱ��܎�:w���k����K'�*����pD��<��s2a�;�\�4�ǌ^�{W%'�΢]ԸjC��e5����6�4M���:4����^߄������O�|ic�RK��
�ԩ��\v^6���JkJ9�|yp%�X�3!;�p����M"���2P��I�	���j���7a��}EEG�����{�d}�#-2��0F�P-��סɮ����o�Ē�i���ܻ f8* ����l�TW�v�-g=����d�h7�Ժd�uG�����)Ij�/�1�^�>���j0,9o�ol�b�������%$��� {���T߀�.�=� G���A8�Q�%>�C��z�0����vVU����s�t��IU?�^��cf@a�I�bw�Yh<�l���,���#mˢ?v��7M&��w�R�.ix��J
nR��(������Y��*v!bJ����� �Žk�Ϋ(����ɮ���3Wڽ?�)��P��В�t��/\5���m� �M_��8E��u�1�
HZ�'{k�r��1Z6���:	Ӓ���9���H��$�p ����`��ͅ~�P�kxO�2�7p[�y�9m���FZMx�w? ��� ��fX�$M����则�%n=$�ifu��<@���Y�It������S'��' �̞,��u���"~���Q����M��@�uC��d��%Jȭ(F���@K��/ϰ��" �R��h2Y����=bt��i|>Q�?Rb_)\��q�HX�e}��V�9��=�<|W8jK�WJFO��=���wY���󻒽ڈՊԸۼ�_�� .��G��%�:
��BPb�1��=O�Qb>I��^_�$a�����B�*�%��5�P���� ;�\��-��m��l���L�g�m�yl�������|�`���j��w�J^NAa
����]Y�?.����\Jg�v_,�4R�Tz���eY4��p_��$�E+�~0ӕS͠9����лsYEL�91�`|n`��6h���a��w�a�+��Z�!c�a�5���ko-�.+�8�C%P9�Y-l��[]F��O�I^{���oE��=���=��#.����M�
6`�>~�����#J�N�_R�yY7n���;��2~���'K3��qN��*u������)G�4�^���_7��z���I��iX2�L��败�6󰓛z���P|�?��=��Ih�s�k�-�3I$�rt��ٹ3�!fbWt��+�@QX������W�
klL������4�����k$�.���T@����5�%�󿠷%��:��9y��O������Y��T������YRT�w�Ц&� A�������nf��Ѵ9*W���>|a`+ۙ���^�p�w������3�?�� �dV'�|Da�В�yN�4ũ��^���7�	�#h�33i�߾�
����o���_�˺/!��ٙ8�0?�,Mw���MN��{���7�B��f��p|���s�(��C���v�$]S��폯���J���+�h�}=�%c=7 �j�;r%�A�N-!+���p���uⱚuC�]s�!i�T���d��ﴪ�HR�×o?iK=Q:�DԖ&/o�D@����l��\�2]�X �'7(�ϱw�_?DOFi�&(>U�ϟ%�5ʗ�l��ګ�,@X<�Պ����j#�hy�w�O>�}8��C��V%���<�p!&fT��fc��-)��d|�� '"������tUDk�7k��G����E!�MP��N2HX]]]xC����P�~}:44�Ɋ��_9�2|�f��M���B.4��l�_�$,�72����Б����Z�Ί����8>{Y�u�
�������8K+����7\� � ,,V�;�y:���^gC���$����a�׾m����O /������Ve���_o��7���}����.���ٳ&������j��/nݺoUT�[DF�^�SQ]=�_@ �+E�[5��0 ��ֲ�3�]-B�Y�fX��@(l2��×�̯$�����_�̨07*��y�g���G�V�\����C����k�'){�>3�-@%-�f��W���7v���$���{��{�y#�51��a����� qS����|ޏ<��D�b@���%�g@Ut篻Tj��� ��KYk����Q55M?}�̤���4n��5���˵�/#h4�$�d3���v#���9e����̛�Y�~��v����j�+�� �͇��y,\�����Z��q�Vgg�6J�(֍�~���J��OJ��=�]��O���]�_�y�V�߶IXX�9Nvw��,�u5��?�d����)G ��[�����YwJ*��89���a������gώONL01���O���^�Z=���鱍����j}�ؾL^|��ӗ�i>�T�V�	&]	��_���%�̌8-#��P�0�{��&yy�����.{�ؗ���%W��b����v��Qa���gy�$tt��'jS����N�f:����.���?(������/����3δ� �g�u'p���� ��D|�y��_�����
h����R�W:l������E^3̋���#�s/�[�>��#���0�;��AeZc��R�֞��ӎ;��yP#lV����%UgX��Ek�t�H��y��iǙ!>C~��n���B�6${m�LF�,��R���]��j2w��,*3�6�S�GmZ�LI�yN�+���#�a��Q�@�r�x8��L�@���E����ٷ���a�pྖI%�p۔+�]`�cY�?7��ͯ��;�ę7"�iߘ"W��xO,�|t}�X�!��=��ä�@��k{D�mS�=�ϯVj��?���􃅦�i=K%�=�y_��	m���xVN��S�D=��k��oz`�Z{|T�l@@�٨�{��֩õ��Y�.UѝS����S*.�Ʊ
-������H;����O�j��_��U�.nx
3h�0�$�ŗ:�?��sw#������v�����5��6��EI7�� �1>K�����N��=>N�mf�JBs����6P���CC>����g�Z�s:���5��{�d����ș�S7����k�Hw�E��)L�������������
��㧆KSt���\���F���{��9=�"���}P� �V��~ġ��:�I+5�a�t���p�~�
Bܾ�)��5��a�Jfq�H�y����6.�&tͶ��Z�!L��~cᑪ��yw�d��A�o�(����z@��rI�CkI�J��& %'0nX�=	�;dx�*��wdj�/礇�VrS2j�?I�F�[�T�Q5�Q��}w�>�1��U�͹G�0�����JUQ�y��ǮX.��9;[֒��:�?�X᜿bk�E7���f��.�y�Z-��b�{/�<��S9]~�2����U����?{YԻg_�p�X]�֘���z�?�m�ֺ_`�^��s��SY 6�±��]�]v���qR��o< y�H�".����C`7�2xL=�0}G�Y����lN!�x��믤e�$�����!�^����������~7%����"�9���fJ�'e�bw����9]�ޣ�O,��]��Umc;����$u��L՟�+���ā�68޴��`�H��)>!ԡK�v�◦@0JSu{Q	�{���J�;�}�;�P�����ÙQᵊ�z�iXt��՝�ϝ��)o���0�>�!񘆆�������Z�z�h�<G/�uu�Bf�cL��>�,i�\K�ұ���'��6��ǖ�-�4�?���lZ�"^�\"��W�1p�A�y��T�,������W&`� �\Y�l��$	FjA Wa�U�p�3��L�|�}я��^�R�?+ş��i��7l��B�������d��4��mw<��{ש��s�ب����J�(�����f������v<�R֖�p����F�bt�v[�ZӴ�uWBG�f���@'.�n��y���N�|���?`���wс��ן����D[a�co�֑��|�������!w3*�O��Aչ�D;����[�3����#G�%fu���^��"�rA����ש�;ү�^��}���D^/MYvo�O�l�й�n��9if9��^�ſ�t��YP7�Qy|ڎ�VZ׎E6��㠻Jj�\j�`��J6Ze2���F
�x�N��-�	�·�>�\����Oa�eY|��B���N�]��J�Y��4�{C��h� ��d�A�e��v��O}՘�����A#O�D���w.s�o癚b�f^�/���9襀]�#�5g�@�H�h��d7��E}�/�DF�#}&Ks��񭭥+mE�w�Mؕ��`�O��rS����1�Ԥ{?���w˔Fl�%���#�i�e� ���Zl�����j�^'{��P2B <o
���@N�������É*��ᨈ�����J��Ph���[��"�Y�� �.ሥf��3¹��.����-rF)x.v���5���`e�?P���n�mdP�==�E��w �6�i��ʧl/���"#8LO�5��6�`E�7�0ۙ!d:�.��^�G#G���=Gq�~��e�
�X귳��R���ՊS�sf�4�,�iӍТ�΋Y�?������Urv:o�彍�l_xR�_l��}[Ͷ@h}[Co�8�̴<Re-ycd�����@�o��ܘ�m�l�M乁����R��)�6���ђ4����h�˶OTa��F9���8YD�H�����D�I����_��n�kn�ٴ�pu�W��xLV	}�Hƽr`����nRNH�ވݶ4�
��ָ���oF�'��L��:��{y��×�9��G�G�+X�'��FM ��x�8m�#T=C�6z�a�2^3�M��B�lXi:U_�#g�
���/�
��df���x�9N�LȂ��<yk�2-�˦b����e��G����M#L�ם�5�Ʀ^jl^�KF���F��ˬ�W�G�S���su7s�%^H��ձ�D�8�|��	��kؓK�XEl��]˚�G��+��	K����K������Zݴ��"Z�d��Ɛ���Ψ8���oF�X4z芭��ܐ��(9{Û�B�}��qw4l��&���4�5o���Η��V���9:��m�|*]$$~)�����s�N"��g��'����<q(���Л�BC�&��{�M����-���[Xې�G
"���)�^,�前 ����7k=�u]��oR^*ɋ쌽�,ΌQ��dc]��\,x���d�@�}W��|��;���Tr�=$�.�v����u�EW�c���AH�9�(,D��?ux��.`�>'��Ǭ����#��2���Q9�[0Z��R��I�?<��8"�cOhPO�6���~�'�s�ɉ��m����'|��Cb1h���'>7����:����?h��p�(���vhH&Y{C]ϟI���]���΀���lL8 �-h�&P�7�DG��5/yvh��Ж���r!@�f���2�mQî~l���M�8��ߌ!�	2�	*z�������|��l���/u�[�ts0vM�r ��"�&���@��ܼ4��d6_q�P��d�@��B.�F� N�D���ק���Q�ݍ�����; q>���V��k�(���1C�~aE�QQz��q�ۗq���۩Ω^49��sS�c��� 椠�j-�b��[o��ʴ�m��g�\���l�q�K,d�ta.ɷv��B�@z��i�B��>�]LD�W��cM a˻�h �"JW��z|q4�g�?uN��Q���T��*)c!M��s��X��>]�6�!���+��Q�5Bv$t��C�pn2�&.=���záMƃ9�W�k���M���_[�_ۼИc�?%e_CdYȀ���'g�>��y�<*��n�7S++����S9��T�%T�����dܕ�[Gp�&��C%��t��]�:�G�&!@��Cܪ �"�>t�d!W�dk�%_�ۃv=���0.2�a!ӠF���|#M0�<�Ĝt��$�K�n��2��|c�G[(�6�';�9�q�y5�,J�_�9�4y�`��!�&��A�3l��Vuz��:d�T���.c���͗�������+���'9�|Ӫ�����M{eeU�j>|8�4	��['�0���_����oƅ�V�&U����M��8��WcH��o�@��G����\ �7�n.��V
��|�NEF?FL^6��K��k�%	�H�(�
�;P��ܞ[0���e^D�)h����w����A�R�8����a��m�*���j��g}b�qϸi)A?گ����ţ_M0�������p�c髙�U:�����$lg���.MC��^D8���1�2Ѻ�I�f�]�UR�1[]YqG�I��u�%8��Y��Ռ��o͏�vƐ�1����tw0��
ht �_�����Ls<JV��u����ZM\�;B�a4�Rҁ!X7���T�<���I�����~� 7'U&T1�8��1�73��Sl��u�N�^�w%���kuUM��=v�K�yh�h�p��Ά��?��Mۄ����X:��n�6�[�156�ɕY�"|��Q88�U��$&il�rӷۢ�5��H*ሂ�F�Hnˑ��\�l����2��Tg�?3��K��ܚr*��LR��2G�*ߞntX(j�7�~�w��}\���X���-;Y������`��"c<tR�3�Wf��֢s�	V8��u��_��e��4��i@O`��&�]]:n�i���4W/z��\��</߸����R��(�߱�lx�T��j�aƢ	�~e�LȍO%���{u?u�I���]Ɩ�c������ߔ������ݜ��(C	'��uw��{��VÝ�q�ӞP��!=��oq�cP�zS�1�,9ǲ�\����f&���~ݞ	t�k9�FJ�0��b}�%�4#��:|�V���E1 UZ��>�k��MT�V��j�AR��g���i��|��P��5ť�z

,�WL���> 5�̗?�߬R�p�=��K:3}fxq ����Ú�.
&s���?�iS��6.�t�*J�=�p�������b�J0�ve���H N^�P�7�;
�K3��c
?��ȩ�2H������-���a�X��g��?w�͇���w��������(ݺ�;�l��53��r�����y����t�2�h�P�0_C���P8���L��*A6�/�f�F�T�Wo΀)u+1fp8NL\�V�G�9i) ����v\�v4�- ��W���0���(��d�*]"w����]Z�5���9��czR��-v�rwuj�C5S޼����1Y]v�rsz�d�����8(:�q���|��WJ1�7�:�T啿�[�{�o��44�,�� �#p�IFO�Q�E�dճ�r����<[��B��d�	�30$����d�X��zL�9n�;��N,��_wT�����=��ob��o>�Y��2_6�6�ڼm��BV܋ ��f��m�s�����'�pB��Z����3�@V'!�M�-ڝ@B�b�^����0��/@a/e-�:��X��M"���S�92U��*~dlQpd�{�:�0���ej���u�|�c	���A&B��FSUG�P9zl��a�`G^���@Y�
8�؃�!(�}r��3�&��I͍���zs5c6�ɦ3�������Z���g��Jq��P���y���2?�i���/C�k�+�K''�1G|U�FoLR@�s=MFE��9����Ӝ�q�)^6�@��.���C��-��3���-lq3���E"��<;���+F>��@���V\��Y��0����p��7�V�lj�qwz8��/��n�_��m�za���6 ��D�,17@���7��}|�k$�5��g'�o'(���YQV.�5y$,�l��bu�k�].�x�|Os�A�Q�K8����A��Ns�{�Kq ֦@P�t��4�d�����^�����r�Z��'�3�'ӏ�
<Q<��E1�i
W��E� ����3�����5�4����� ��� �
�g_�t(��3��f�m�����a�^��u����c�:�l�=��߽�k�x��w�pƓh�f����@��v撕:^2��q�!Ɛ��2��a!µ��yO"����W!)����'��s�Ut�����ț��g��0���;�|EA��Eoy��if��hq��3��tk�0�����1��u8�(wi�C -��<��c���A��Y z�0�#�cӍ3��>���t�L�F���?�:��U�Ze�,%\�Ԏ�͑.�H�~����f�??k>%���_��	��,���K��i�w���@��!e�Ќ{��J�_�������mRٰ��#���.
$��X����i�x����E�>�Ӿ��x�H�+����0����BR������
S�@�����'� O���+TQ��Ø8��T7�<&� YAmB���y�*�����������Ic�\ppc��r�'`�D=��Ӟ���y2���Ց��g48�����K�*�9ybA �+��b���/��!��<k�|�պ����&��%p�|϶�Y��w�j[6=O�\r^��]��#i
�+���O�ۡ���?Ì6b��d(S�i�..l���)���}4(��P`!31�H�c1��y�)\`DL�L�����LKUa�H��yC��3^��o�F������c�D7� `�����6�r6S��]n?8Q�P#��I;ľ$�/��:d�˗�UN+1�N����X�:Bg�v�����msV���O���m��v$�<a�>9�[����8�I� m���=��	DSV�]3P��9�uD�4�(�����Px4n���5��w~˯8KES���e�1��T��O�n�9�p����:RtS�@����w�i�w�7���Fv��� �u��|=N�ٿ�Ƀ�=j�E$)�7�8uw�&���e���q�)e�@,$��V�n��͓�!ǾM��G��t�F��\�pE���_���b��d9��uZ�0�>9��<�WX]�?�K�D{W��VW�v�Z�`����)�Nf�®��7�{��˜���{�3jp��5���`����z)I����T<�qf�
��w��|�mw�<Fk@�7, ��îl�O�6\8n%��d`Ny�j�� RT�P!�WR㻦�o����K8ȭ}�	��\�uS�_�����Gm���n&���T^K(`�l�c��_S������d6b��F�n�@F~R�50�vW��AB
ԍ���ۂq��ɷX�o���Ft�U�w"?�or�5��:��׷`~� �`��o��6��&I\�S�A�����0!����ݞ��0geh�pT��w@]qp�	��8�S�*�:��g����1�u����&�JH^<���_j	�ѣ\��_�	a���t_ ���"����n��L�ڊ�rB�� �É�3GB�%@3ϸ��8l�x�{��@�=��F��9�
9�b�����@�-�s5?�<J�c���!Q�f ��i�,�2�E��{k:Ku2扎2�m�/&OI�,u�2�n�!��
g��y�>n��π(�h��e��_0i���G!���uk��R���[����N�]�8T��緟�QA@"7��ư��'�{�\ެM3�X���B.]��%`��A�����Op'ջ��8{��\��h���Yao�t�aW����m��WYw����]	��%*���/\����f���`"��,�aY��,wnm�]:��g�ʷ��q1��΄AeF�o��|�:�pg>�t�[�3I����MX���ʓ�p�x��YS��kL��_�kPf�x�<3˜kKKe���y�8��:�P�n��|8X$=-8ʬL���*��A^����\�{�'p#�
��J%��Mse�v�����̰��I�Ɠ���F��ڪiH�Y������&���e�*�v�x�����l�D�q������/Y~xw�m����plv:sjz���$rx�����d�'�gLh�8pcǃ5���㔛}N.��q��q��a�fX|{�0���mt�a�H}�Ӵo�r�Y�r׎�����X�)]��8An4�D�����n�����⬫暟���Ȋ����W�4^�O\rLNV(9�#w��Lݾ$̣a�!��!��E����D�����Qh��4Ç�&�x�Vxsh��Y��e��/`Ws�"1��aNW�0 ̤0Ͷ���8�?	
�tq~9�VR11����r��>Y����m~-�I��<�z����_�k��{�k�Gpb\���'����c��?~LH�9 1'�55�IKTw7��F�z)��~�>������Ж�=�Ҿ���ny,Gf��[�(��n��_��� ��T�� ��&�+,�Y�,�c��j����r|3w��x>�j�������H��q ���Y�
��MA�7C���:::�Z9����޵WC p����`�[��i._(G�vG����7�wG�농�ĎJ��`����������l�2�*��zX,XXX\��GB�X˘Dv�EvE<�t�'���%;�b1��"��YFg$"N����ب��y���W���.yf��?������1O~��aֻ8yx���9HD�l���_�?sY�k��OlO�<Z��a�U[�>�SQCbbbҸ�Y�l��\�s��a۟��0�Gke��2��h�׏s����,s���@tΦD���z��z��E産�t���#.�E���� �,ݿ���p��X���W��,ⶐװJ�B�3�W6;;{|����m��C�~ZZZ�L�Rb��;l�滻���
�����o��X$+ݴv�\��މ��{����@�%赛�����}��j��ՀK�ǖ��Ѓ�q�9%�3o>g�U��L�Vϒ��mW��O��cH�6����ډ�u���.3	>w�j(^k���s���<����9����QV~Bbs`���#�}�i�����=$�Օ��ڹ#�� �v�~���v[s5hD�������x�l|���P�ӧO�۵B���������57?�'I�f(~�>\'H�cN����}$>ߢ����Nd9XT:E����5�c�:J�BW�<9�����م_SܹM��q�����FFI�/� ]�c�G�1��K�:����L����B��{bv�#ㄸ]�%t;� �P%㫳
^��a�p�m�2���s�Ή��^�vi��[���)T�epp$l>��r��+[��s�v���4+�1��V��1�M�iZ����pq����鮮.N��<�Ł��x�i��$���2>i������ ��q������f-�I��r�����M����Qt娌��~!4�}����Q���e�]��}����f�`be�H!遲���ߌ��S�m��_��.�ϑ��|�#;�K�l _��5�jY_e���E0,$Bx-��u��\q�=�Nl�?� x��B����l�������W�Y���I���JK�L�Go�n�VŴ�8��L�j#Fw�U]x�)I�ʭKG҄��u�t�^s�t�jhnRyy�����ɝ��U� ۟��L?#�h֑(�_bkHAI	�����:T]/23�,c��H�ɕ�B��V�'E�k����Xcz�'�����E�ۉ���=���4��E���9�����򠠠 �wT�uT����c��{'7�swvgN�:����Şb�K�9�;}ee�x��/_��k�F�a��8��e����s�CwX�a����������;��$���
��)�Άl��aέ�pt4n���:%z���|�U]N��w��גۨ��Qv\��2i1T�G�Vjw����r��yb�JɁ�^T��XM^ja!w4�����Z�G}>R80dt�&�ݭP���N����:�X@Spc��$^w����ӘGz��c���b�Gph�L��t��;�[$���>fN}-�ăik�ͺ��"P[w�W��d���`�F���i�i��V4�o��w��� TMMM�~�V,������3��X�rkR�vW�s'ܫt��/��Y�*�Tnh
	�q�TQ:�����P�3�מp�Q�$AC�[%�#bâ]4�9'bm|�
�UH�Whis��(y,��RN��3�Y�J'�طq���=������f^�dp��Dm�HjU�����#�$�@T|Z���y,�og"x�#�ӡwd��k��}����)�I�EN3@m����̜��Z�[�/)�J����q�,��Xa{��
������ҍ^���M�/ȧd�w��v�����x�������Nw�p�]� �f^��Ǻp[y�C�xl�p�OTtql��A�����b8S���K�z��K��|��#���i�����^�X$	��+���A�ߝ'Hм���W��{+�*���1�^<�\�(�Ъ���a^�͏_���=37	������Y��OB��嵫P�*����h�x
Ҽ<�d�^��^}V��ӷ�A8,22R�e�d���|d�j��aܵ�h~nnu%�Kp5�)?��@IQ�,>�`d��9��}�.��8�� �e	/�S6����ݳ7<h]-D���@^W��sqA���m�°T�r�m�855U�Ό|;7�!��ڦ�p;�ջ�pE?�ԋs@ڴ@v��,�e��i4Fܚ�^��Z�k��՘M"�R�hUnߣ��c���g|$獭���������|t�x�t	��t�*�M��]�5�����i����*~Gǔog��g�d�EM̱g�  �v�ݪ���ٌ�ʍhW{Bυ���GUl)���@���/|�'�ːe���:^�����o��c`b0�LCƦ��@�@����c��cB�5v\k�H\����$e��M-Q�J=��	=u�p��"k�"ʍ�G������4O�����5у�lJ�c�v�m�f܎�݁�m�#���uWt{� ��������s271���pb)))`b������R� ��M9��W&���������l8>�b� "�@��M��n�6�&�]Kb�`l�N�oۄ1�Ekȍ�^����C���"�Q��^��Ғ��i�X��n`�b/t��0o�R��?n&Ђ��Н�{�_@2�Jr#���ݷo��|�������ɵ_nɄ����g�Of=��S��˴X1�U�ck�C�Q1\�<e�_;���^�5F��>*?;/�$��Jl�]-[+.�Yj�������{���+TO_&xƈ�~i��0�b�YdMdz.3��F��q����} X~G�)�'Lt "�bW��E��ҟ�P�&wpp0���]���-��%�����hN ]N�A^Hv[�ܩ�z�P��h�%@�����OT��+�BE��2_�a���(Q*Q;��;a�I�`���v;O.�gR�kC�x#�2Q���K�~2*�5����^r�Z,���;p��D�8u���� �M��>O������z#̵���� ��T��.�%�����>�G�5\`G}�.��"���[��0d��3k�1������,�\C��r4V3++V�'����h����I,_�\�0�����Z�ͬ��_	�Fjt���SJ��O�=L�X����_V�]Y��%���EO�aǞ6Ԛ�ǣ�\*s�d,�����f)��-��×h�,@L�ХE/�#����8;��uP�$Q�-�Fq�lnZ��������W���RT����B�MC��6�**I�?��ZXV0K^"���<;Q�(y�fS�i�Z}�D*�ʠhyJ��?|���B�
������ ��E/!iH��N=����)��^R�T��,;�H9Ȝ�i�_C��{���J��f�����#���'����Tם��!ͤ�a��C1ϝ��;{=�7\�PX@��}w�~��z�xd��c���n���.�k|�sKH�V�%�p�@LM
|OZ��Q~	`��0m��լ�87V�|5���t"�;���G��R{Ǡ��oH��	��եu��l5�J�bn�M�1��2ۘ�w?�J��ݏ�>�0�Q�^�%�w��X���ݷ�0�?���1**J�43�
.lU�XӦSl�c���-�SAج�m4�}¨�f	a�HN����|��Fc* ��|�.A()+�XJg3����Ks��7UZ�m�.b��2?���:����XXX�;��q^9E�.v��ʣ
`���!Lllȝ+벧Qt�S����#w7����?�@]��z�'���B?��=�!��,!�	>Mש����齈�(c_<����
E��ýG�n^�_hXzCt�������̷�8q��1b�Dי�'����?X�[����a���=�m7V���N�C�rss��p��B';i�G�Z�Q�L���U��^_�cV �|ϸ]C��wj�v��G�H�!�7Vr�F�E�G��5��]����7�E(�{��� �Σӟ�n�� ��8����yN��W�V��������k��)�l*�ţ��eL��=d�4,������N6�D��\�ӈ���u ��ƭ�̈O�?��ၭ-��k��jzs�\�Ǻ���M��-���6��k� `�.0T��s:z���@IQO�&44�7~�7�1��V��j�m��K�z����oݻ�i��r{o@�d O���^V{��}(&L�{3�x����G���� �6�*A���i��
�19Q<�ZC^�p�(S�ۂ��n-������|��R�f<�!A+'p��^�o�:���[@��=-v�h��u�H��F�&U��T=�N̽����,��4�IwI�d�
�^426��2�.�Z6i;=7^咽DM�Z�T2�dk�px�'�@�'�YK��T�"��5�˝,׮�:������D��
��?ϰ4#uNk�N�Dο~%�W'�P_�f0~4������P�Q�v"ĥK����}����� ���ڵ������#qmƤB�A������r��^�y?mP��*XU5S��?�P[y0� ���t�IL��9o<o��M�%��HP}c
5,���2��x:v����%P4��1���˯�Q�^;k/���3¿Vп�I���73=]��m~!�D�&�΢Jo�_�	sΉ4/�?ox"��^⍯P�jj �b#9^�X�v�JW��_��xK�s�am�K_)ƗS��^�w�L����֯m���[*2mbV�����p0�'(�~d�W��\�$�uШ�1~.P�}��ff�߳�S L��@X�_C�5�<�W\F�)?��������D[o)y��|'u4������n�k�*��(���c�ySʢjq�q�9�yl��ĳ�mU����/���hc�Ƿ݇�`ܢ$��^`����1qG�kׅo�^�E�h��@>�d�z��ݨ}���J�j����wr�<�>�#QMYlݫ�f�_��vR��.+�6yE�u2�25��I-Z�5���y������'�����u_��%W�]�N�,<���C�3���s��|k'��O�A;��+;���������μ�2�Z|uƫ��+z���8�`�����3{=�� �I8�a�[�>^ڎ8O���M����2�`R/�����9�I�HY�n1�\*@���vuZ�L(�E$:�`�x%�W�GS~/v�͜ ^vm�h��ƍ:)��L�\��O�[_��
L�}p�Yi���C0���
��k�ɧ�D-z�u:]���L��O
.�,����>���������8��(m���k ��1=}hBK�ӎY7o��f!�.[i��)�A������rt)���}�|����h nc��Y>|�]#{�x]o_�n����~� ���v�-x&�D���gԸJ�oϩ4y�as����N���ɠr�L����e�/=͎�	�oDv���ّ��k?��܇�5]�=
k�l	�Q�XX��]+�+�F����yȁ;����Н'�>LT遏(�0��TJ8aH���9� JBC��Q?���b{��+[�-�š���d[^5�f�s�?����b��9�܁#]���!On���nwǻ��9l����,o�.�>}w0��_���Ł��n5�C��ybv����,��F7���=<�9��}�뺝H�A�N���`4Uuu�jO̅�j㶨Ɓq��1�e�� Z�`F�}�Ҿ?lU���~w����'=f>w��2��x2�D�����B��
�l�m���#/|�O�w*�'!Ѳ�zd�6��J����o&��-���@#s�
�C{�n'�@N��S���i-�L���ȵ�M��}
��׼���(ľ��,��0�{���0 "�UD�D��̳dH�NTm[y�� Һ}$@�C�KG
'����n���i�.R`��`_R�zXM����8��������"�b|q��ദ��4� s����F�ڨ���A�mN7v�E����K�&J��ag侴�ueF���O�	Td^?�����/���>\���q��>�p�h���.�'�9=�����Q�omĖDN�֘�s1�8��P�J}r�s�v�����I�������L�c�����u�W�.iXy�1�+��M�0�Z5����c9�R�54�<e~�β�;�Ґ%�	W~zg��7�(�.Um���^l@lQ�8��'�t����/>���r_�~��Dӻ֛�V�͸7�i:����ً�2�ʦ�5��z���;�[e��,�U<��l#Ǘ�&j�E���Vz�R�1�Z�E�ͺH�q�}�b��p���T��'Hh��R������1�L����/~2S-[�A����ݽ�Nse��Q���+�'�6�^'(���з	xu�����9ר����n����F�'��T�i)Ǹ�	)ȩJ��!�޶��ab]eǭk>�`ڕ"njj:��g� ٽ7����<O�(�z��j�������>��HO2��7M�s,���,�	�I�}@��!�SIW��p�.�
M�q&b�nFù������&���~w��5l���)��`�c�M�S�o|��ds�R��u�~��	g]\��p���x����gU����J}��������	)lT���Ue��8HH�ֹ�X�W�������������}�N�6J_h���5�Ƶ�[�N��� tz�պ���PUU��ifn>�(�#E�\�'{BԹ���yG�~̫c��%�����С�4�O����2���$K�j�U�b�:$j���;�c-z����4�`qp�l�ݘ���ǾbR�>\��6H::;wV�455u\g�W���&��)���:�₯�A�!�OF#r��-܈\9��Rɬ��?ʾ:*��^P�c�@@�[���F��.��N��N�.�����;���{���}�}k�Z��{���~���9'����[>��K��R�
�7�R�{ɚ��pW�=�7kV����pe�����O1a4��yD"x�xY�ևih�'��b���-�C��� �Z���)��+~<9������N��6�c���3�o(���..��8�<.�诏9���j��?��H2�SST1;_b@E������y4���v�U��M=�QV��!�F1����V�����t\���=I�����(.�r�4���]���xiw�螟�%W��gH�?�~�;��ˉ#l���bY��H��
fm�=���t�~�X-������x�+Im����|�}�A���I36�F�y�`��
�J�Vܝ?�Չ$���yH�Eu�Ҁ��|����Z
>ĥ�	����Ӆ�#3��^�X�K�D�,!���WFqo�}zi�8^f���{��!L�Aco{F#��6@���=����a�DFu��m�n�9��XT�R�k����dE��?�D��<�T��X�=~���� �&>�r��L ��JB ������l*�8���]��~��Dk"~g[���w��8Ƚ�E�:�l��5~��68�#���C 9��䫴4㔯I��w~x�S�y�zF`o~i,���	}���	����'2f����}�py��΢#0�|��9r�맃0�x�]����(�s��)T�������
T@�{T�k�G���=�⧮�	�1�L��~��F���bki���s�����;ӹ�;--������y�MU�&&�N��K>�/�ͼF��`��bP]z�),n��1˦3�PL��������X����v��g�$ɝ ���K�v�oo+LQ��>�6����D>;��Q�W5��O�����Q���.C<N�%uKf�YG��I9l�_P�ݻ���Pb2�ǵU���NwjoW僕���nr�+V�{r
�b����q,��c�aRo\�_i�}�=IR��}򾡥�ݘ����e�ͳ�p�zʩP��׽t
�N�C��b~?11��q�tņ�Av�����D��`������I�f	n��B���(����49�!�����[���mQ�]ulz[iAH��s����mx�rh��h��Iw�U�9�0{8s�됖�n���X$|>��р׻�i�����V���$�-�h-w����lt78�B�	��{߳�qG�,BED;:��s��.P���߬��G����D��ݵ�v�s.\�GMș/D��azq!����-�ta�k��"�2�t��q�*/gs����yo8�Ӂ�Ũ$M��}'A\0��A�U��[�gjͱ��������oÁ빧_V󢃼ff6'�����U�ƣ��K�h�J۶��`d;��@v�1��q!b�h����xY��d1��;�y�[ M*�������x��L�8�2�GR�䎳�cx,���(���h���/u�� Y���H�k?a^U�� ]8Z	��Z�H��v��3�ǭ�
,��6�+�	.��dt:[%i��\�l=is �_��8:�32��V'�XQ���ӤN�tq7���sK����ċ�ۉ#@^^\d�w��A�?:qվo�256�+��h<^�'��<� ���ZA@z߸��0�v�a���b�Ӡ�[c���H
.HD��7��c��GաҜSxP
���L�/o���ޕ�����q����>ɼGR�ᴴ��U���/ͺ�OU&i��oog�cIR������[]����� ��������/�y���P�8���Rd�[��uk�?eg���a���h� +ڍ�	vW������ގ�9��d�β��fh�ֹ�]y�a�J<V���A'̩N	� )5�v��ao��ս�*u)A/\��5~�-�0(\?}�j�ύ�����P!7KH���4 �r��tooo��o���;K�� e D���?��B,�kd?g�ڈ�ѽ��-�+����Se�ZtKw�<��/��������@�@�մ�J;@N�/�Q��S��h��MCAR�l�  �*���9]�l�\��LCI�*􊖖�_�~�9�hۤ����]�6PN�Q��A�%����IR���g��x2	���X��/I���d���A�
呪�ת�P��(��
Y��~�ID>d��x����I$+I.x��*-��� z�U\��B-<;�������x1<���A$�@�)IŲ>�;E[��7U��G��΋qg�ʇ�\�*�����/��:���n����۪�s�9��X`Tm=�3db;EZ����hMSX�4/:�h�F5�J�Q5#� �_����^^���"��3C��*�8�SR��A[�1�k�Ӎ.-���CU�,$<[Kz~�s��Pr��&��sV��;5.�z��JG�uwu�7l�Y�^�����\O(o����hD'�P�Hb8Vl'm�b�m�<}��Ư�;/�ʜ(�k<PH��6Z璻z���7JN���?
X�O#��{��~���.�~����\�����oGNm�s"�B��8��Hnt0�R�gV�6�-�vB�����-�̫�8..��E�X��p�`����Fn �w�ޞ�KPq� /���E�����}�ţǫ�{�A��z�K�ޢ������C���80���8^����7� �8b�N�+e>�ď@�f��XB�GEK%�����`����C��W��k�o�6?M/j�]�ԡO)O��hL���t�R�����x�P�w��l�P�	�?!h��'���y;�LMM,=N&�?�3-��7���.mD�W�N��3$��Ƌ�{���p���j�-^R\�<�EY�|�6YM���eGǷ�l8�����D/P�LD����a5�<	��>�M�U���L-�D�n^�Ի�ܼ���A����

�y��{�K`�H�8`�L�3|j�C��K"V:��Ǿz���Z"ל��h����6Y+-eVF9+�üb�b����}����B���Zi�.�HIK�ԗ���f@�숞���5��a�j\?Z��ɩ׀��0pXo�s���[A�R�m�D��?��ҁ�K��3��Ӑi�T���'X�PQm�O�NW���(���pX�uGP�	U�;�#yJV;��Ў ҡ� ����Gs3@zy�� ���o���v�M&"2�� ;=�](�	����B��9��A�V���Ư����68*W\<�[u]|�Z��n���l�>$"��7ع>N%�8�X?����{�S]��;��w�;i�a_�FY8���ZYI�U{��/�OlxvA���Y����E�.�>�Sæ��X����A��M"�a��o&V���7	p����!��}j(T��ߞZ��K5��:k͡�\~���7
-8Q�d%���& �P�r!���K��O�����#;Dl�6��M�#!TƐ
�/�K��3 ��h{�f��v莟wq��<�t/t�D���l�����1c+��e)t��4L�>xLr �n�t4����:�.aY�oG�7�\��<���o�_�nOO�߄.������d����-	C5`�a����4��j$jΦ{�g	��*0�;e�yI=�BTH�wf�����޵�s l��Q�
�׾(8K�σ�S�$y�t�ϭAx���d����a�'ՠ'Q~\}����ka��~%zЎ6?ܡ���#.�$��g �@|2RE���#p�lY>d���[Ծȶ	�1X�r��W�ջ ȨC�[$S���;�SSfn�*xP�Pd� �|»"l�NAϫ��O��+����Tb�dS^��<,����~�=�à��à�@�[ݻ��?#{X�FU�s+���>����o��/�vi8L�c�2� 4���U�9jcT��&�Í&'�@u]�!ujE;(p���FaU��8���X�6 �k��C7�b5/�-&!7�~S�"l�����\#��7k�B����I���5�0ĩ�d>#����3-�dL���1�S<|�r�V�ͳt,��b~f�FM{غ�Vp1!���`W���7��Bg���w���R����-��x{L��/���`���fš]�5�k%�&���ˠ/)qh\�}�� �VCҜ�)���X �4	ؕ�}�޺�X;��T����_�ᯉ�����H�M��e��P���Ο4i>�ᨺj�	���s-��̓zL2.fW|Ff��˶���8��|g��A`M�� S^q�FY/ݥ���^�Y	�>���L+��%O���w�	�4v۾xsF����َ��HZh��6����A9h��?����w�P+���3�z�"����ݵA 9Z �E��p&�Q���f���#�u�j9�!��+����A��ܫ��<���� ��q~

$ҁ7E�l��%��fCn���A�̰/ �L%Ǡ,)�)�4��i���MH ����9�V_�\�x�9���. %8ںpa?��R�2�n�2�&p������g  ��x��I�� ���"w"֏�O]�Z��U�< �uJI�VN#B�8v�����������d5X"QTV�w�Lp�@'i�)�[�>|��`>cuh����ŵ��#'7�o𓗃�� |5)O��Ld�d�2 �/�Qs8� P�@P�d�p��a`�g����j��>I��^��W�.l���KYi�V�p���ǧ����b��$IMyz}a^^ޘ���h�hQ9�~��71��i��~oޘ��x�	,�������
�^����1B%=�4��'s6F�b�\� �bl���� ���>z�0�2LϐP9�1�-�Hb��P`<�;���,�w�Kp3P$ƅZM_��+#��,�^�������`D�t9�N��N:���������{��%6��N�d�&���AsXjt[�rԌ�&A�n�C����r�U80��F+� �q��猫�W«�'��J���B��[ �{���@Lu��������"�	���b��t��	����T�d%E�6 ���O_V��>M��7| c c�O��
2w���}��@�����jO������T�~!�Fc�U���kEܘ-��@�	ďd5��q�� 0��� ��>1qI��N�	���4��@e��V��%���``c\�������#���'88%;�@�AK���#�n4���.���f�~�����\:�5��iL�ڕ���I�
�������-�������Z���A	�f��V�'啛����� ��3S�~Aq 7-���~ e0H���5���*V�6ߣ��2��t�L��$�A���Rf�ƹH�O�nG&oe+-��'wf�:����{�.��)Y~�b�݃��>'k��������5����QLZIeN�*��Ta ���^n$���ട������Ӄ��i�M�u�њ��3�@���X�٧� � \��\�9�m �p��yW:M� �G�V+keƒB��[��J�^k��s����bj�Q��py%���i���gacի��POE��̠������r6�n���6�n���i:-E1�`왿me�	@�����	�\�� �*�i��o��,bV�$�ܩ��~�k�p����aF��L#��@���E��@n����T���`#���ģ��,�Z;L�O`@0�Ouڷ:㧛���
X�fq�_�R�Lu����dHQ a%=-�i�M�l29��'a�]��$gZr��P2�VZZ������>.* ?:s�N C�/h��ZM��8�Ef7,�������z�(�Q&d�c:��I�x�j�(Ꞿ�w�
�mh�����1��C��7�/4O����R����.�&&�wM��e
\g}�%6�CT��`"fm�^C-�����ۊ�K)X�yo���A�8k�� �8�E�PHKo%�ؒ~���&�f��� 0��Ɠ-�"%��dff� ��IDʡ��zzz �Z��tһ0Ǚծ1��1���D��s�{��-d.I�8 ;�_	��w��\m�x<�79waV�Ţ�H�ck�k��0e*���4-� ��h��tHC���U�hύ1Ў��, �C���#h�5�����``���w!Ц:k�̑��(��޼�,`���2."�?�� ��,z�U��N�R�Q�<��د=?^�sv�6�e�uRR�U<9�Q��ičLO��h:���~������߆�Z�����"�}��KQ�����2���@Е�}�C�@cjb��##ZM���z����c��y=��T6%j�E�Π�b��������gq�%���������{Xb�6ȵ��>f\O��� �`�Ӯ����z>�4�W��"��ȱ������ı�=C�k�߱/�	�".�SKJXz��AV�\�Bg����e��ӫW�#|c��� ���b'�>N��c�D�'|���B����G�GV$��#�b&�	����+�Ʃ�K��C2777�����ܘ����_癞ӆ��#��	SFGG����D^N%h���ʅ�6���E5�q4��2�2& �hj5`j�q:�4�r�������������(({41K���M��k<CXRs4�~pAT��q��nC[�������ʅ��#�� �����+Eīz���9���w�3 �ϣB:���H@�H@�9`3Tޘ�;�6�ZL��Ow�%�܇ ��a����M����M=��7�����x4��D���2����J������B$©D޿�z��5�uq����_��e�c@���t���D�dL$�J�����cs��?�@@�f���E�g8e��| �Է�
�̮�Mޠa���Ke�|���X	ҋ��	������Lǒ����?~��L�l���`S�V�QL̘sJ�d���t�� ���$���y	]Z��� ����y�Y�[hӠ0�Y]�����6��y��_	&ڽo�^��y�_ɩ��KF)������<����+��JE����L4����c���<�F���{n]�iJ����;�ED�8�i��Ñ(A � �W.�=0��\����s�Ü�ZI���FD��g}��Z6�j���|�]!�q��&~5����SDX�c��\��~��b���8'�Z���J������7��A:�%�c��[�yJq�,��&�M�5�G�3 ��S�r=���9E4��
�l���C��8����j=i��s�o:���1L]���V;l�wgA.ic
�zy=e@]{��c�)s!�H�L��m��������μ�(����W���&��_��=��ޘ�!�ٮ�ɯ�H��S������{2�m^�Zɋ꥖H�OS����3ӬE�������	��{GdA�"�7Ƞ�F��F��?�f/�x���_~���;*-�X�|Ҫ7s�'�{��f����z�Fڷ�N��TС��][F��a��~��Y�`���]/{�`�A�?/��0�~LmaڵBW(���k�����UeX۸�N�c:��p���2�^.�ذy)p�pnu����v�WO����o�]8��x� �⨴}#� F_d����,^�b��g��q��l���P!u|�z�b�!��~͞�W�o�����l�,��'RS i�߼SX�O*�\�&Y�ޮp�t���q𒔔�O��(�%O�i�<�5֐�����h[�7��1@�y��((��-=a��bŦ��խ'.m,cM`8�'\�+�/bu�`j�ze�UW�]H1M��%���ȃ������U΅���"��'�1����#��6�ye}!)�^Z�������â��A���i�����p��X�W[J�OM���	��f��]D��yV�|�T�����(�!�镞�9k�T�ǴRri�џ6�Qp�����W	(fm: �K�1|�W�7yRn��.�K�8u�<L/3]:p�$Y�i��T�`0O���B�%ý�k`̣��t�[�1����~b\�����m�jU	�j���̔O�;��&`f
���ꁁ9�Z+.�ԟ!;4���?!8�#�@�A�(�}/�j�r������Ɯ�,d�=Q�@�?6v�6�*�&+\�.Y}����k�Zί����8'fL�1l9C�N앶m��L��Z�]V< ��v���.����oRT��	V�dVm8@�Z��0��hȧ�
�R���I�=݇Z��9�Loy�_���OFd���[K`6:|ۏd��^��cvb#�w�5�*&2z��_����
.�#�'�@	g�P�Ӱ�|���ڪ,�spL�G����u�����6%���j��<e���B	GN��VdZM��;%����'�޶�d"��ģ����\��LPKr��5P4]���=��w;��Y�]럏��@rWj͋�OS*���O5g��m�_v�+���'��eny�AA� �,N�`=��Q6e������r8HSꏒb�7�oWh5�s��z���1[��+������Qҥ���|��+�}lB�p��z�����(!\�˖D�[ה��f/�
T�z��f=#�Z��j�pq�,D4(��p5ڼ�t���|��L	|!n'8���r>?�����A5��F�6���ťK�b<�ItG��A�j�����Rp�&����S��ت28u:6��J�
�[���<�mL���*j9�@D�:��po��2 ^��3b��� ��L<��;ӛ��/����4�L��)�k��k���!y�*���%�ɑ����^z��
W�Tᵏ�!um���w�8�jkK�cL*Ρ��*t��C����ccw��K�G�#c��/�>K	&�g��Cv���j�?�-��N:������tmv��zh��i����f��\��~~�qj�ᙦ}E�܁�ɏIA�_�8|��(�X�qk��N�+�f�P�yY���i<r�.�����&�o<}]����G� _�������Z�0��D"�>҄%��-�
&˭2��2��UE�"I�v��*T�D�\�h@�ݙ�JSuK��:�y����"����'P��7�M�iɤc"*wp�9�@{�~�mf�c��3N�Ze6��𯯇��<�1*ac�c~J�Sux{��kNzMԹfa\Y�	����ڏ�Q>��_�B�Aʹ�����5"��t,#6oS�CS_>sJ�9R	����	�%�k��=!�M�о��N�޴�:�nrr��V:�E5�!��1��7v��k��H���d)&�o39ݞ3z-�&R�Ѩ&�S�TBH�>�����V���mI��䍈��{�3���b7�8�uϔ�����F�sCmE�������ő�-��L!��Qb���#R7��C��&5nx��v��Z�â��kr�a"�`ơ��OFm���B�h��k�_�&�6�����~��r;�m����W\?���0��xም��i��Ӓo��ɍ���IS��i!�*���PV~R�JܕE{��M�:�O�#r�t��3a(�l�C��w�Z�>,`���`�gs�w[�������\����=���L4T�l<��b�������w&����1��:��qf�ЙC�xgfz������GG��%s�=�Vp���]����ckWW�t���o�Ml�+���>��(��m����b�j-o�+"|�QhF���/D91�=�1��VO���5M�{���{YH3�&\	!�����`���q��\���9��8; ��^���p؞H��j�;Zv��n�����.��Aa{�1�q�SF�m����c�Z�Oڠ�]3���U��>��p�ٝ�ug�ȪF�[�!�= � 9��PX^2}�%����D"���tul�����B�owKn�(�-���6H���9P��P�M��Xu�`l��7��凮�6�`*��g=�V��*��ay�ݎ��YR]�`ƫc��{�4?!���7��IxB���!��WC�mP�7-��f󿧕���9�KI,��j�u�L�
~�v��n��:��d�u 	��+�h}�?y�qg�__G�FѾ�@Ӫ���2��l_���2s�VbŎő�������$���ݽ�����&�����=�Z�c�o3�ZH�?JG�/0�?Xxb=''2z�wnsk��]���@�it��,�η��RWo�\2n��vq2�"ԌY�	�x�4u��ac@�b���[֝�AN��|���zn0F�S�V��+G�Z	l���˅I��17�R���e�勳�tH�{E��#b��8Α�*�����B�U�|u�h+����w~���������mGN0U�~����.��ʔ�2�7`�CY�$DD��ɵ�����n��G{ү��$��>3�N^�e'}/����p���wo�7��7�·^�-N �p%SAWڭ��俖�)�trσiyhЩ������{���k� ��>s%����?"0��Ƃ������G�i{�gv̇}�59����6tm��)ũ��:�m�pw�'_-�Xߕ9AF�]���5�מ�N���|}t�]�F��u2�}��*����<��0n'J@�ȉ��5gJWe�~ܨ	jH�<2®�����/�:�i7���x��m;�p}�	�U��E��|�ؒ󀑢Ì[�V�c�R��*��
u����2�~b��*�m�qQ��Q߉̚�l�`l���&�2���+�?-�1�/,�"���.Zo8���4?	=�����&�K�J<(ެ�xH��-�G�nc&:���Zؚ��Y��99���e���]�ځ=Cv0�� �Z#�"��m�mx�4���K0~��8i�S��>[*aO�JmH�;�}]5�ӌ�E�nHL��0��<�F�W]�9��z����!2⏱���s��JXH*�ۇ<	��Is6Woj��-�q�8��R�R�Ȗ���21q��#ǖ�����c˻����XXV��ٮ�����;��XN��$�͚;�-��U��X�Ol�-��<�2��3m�Fa.i-�3��^h�xO��K����z�/~����35gǖ!v�fqJs#��4��^�<r�Oj���o��
�ƍ�&Z�~X4�+�N�u���z@���K���N<9���\�?"k�38d%Mv��U���T�bg.��m��W������9âmE"e[lƢ�):�IX,;�g����d�Y-uy��V+WV��W6n{��8��:U+,,�E��W�m(wߙM���x����{RpR쳪p�p�Wr^6�lH\1�g�fƲ	9i��0��g|�fłԕ�g��?�r�U����@lǂ(��W˓�b�{[���C�1��W��Xj�D��Y���d36�Z��ڪ�3�Q�\�3s0D~n$3�v�>�QQ����怊,r�*=��q��]i�$%��k�)}6+�B'�#�PV<>��|��-ru�Yr�7�b�����n5�F-ֈ>���*�����V��F��m�GT���>����~���� �w��#r�r�k���^<g?N�D9�ؙ� G)����C\0��ؖ6���ki��fbFk�M*���D��8=}���Bn����՝V�H}6�P���,jרD����h�~���gu-�LE��%������08ߙ�Ht�k��M��=���HyIٱ� ��RHrH�[ t� �k����;���4խd�U��Aҟ,ז���b��G|�z�n/oߎ)xFJ-�r"B�O�3fe�:-vp|;Nd �8CIDk�k�k/2\�vb%��n00֘�+6D<�$�9��%�b���Dn�7��8T3��Σ�9��x������+���QO�O
�,�]xT;��+�a�]����ϵ���tC���!��8B$�����2#��o���,��lI]��0���Nn�dpj�F�R��(�O���ď�{���)>]���S۰�J���f_��,-���T����3���[�G	�� 7�^���v~��X�"4�,k�������`��@eT���M�#'.<?���k��N�oZ ���G.��1�b� ��j�c5�L
�v�o�Ww4�1W�#�5<���Yk�8������,��d�E������V�]�#g�e_Ѫ~�rti:�*�aT~Z�:Ms�|��`cb�`�h���}�������Ǉ$�O��B��S��uV-^�M~[ؠc�'����3[�l���;��	ɋ�vad���u?�-kb��S�jq�~[T����� ���4�p8-Y㖐��;���.@�ɲ��RT�t�\���/���4,�@�����]���D�%Q�^X�S�|w�E�����)�����EJD������^��}��|�!��Isz3G�W'����
�V�^T	�+��J߄��{bb!���y�3�@�$����������c�`���A�x��!���8��Ǩ�ݲV�&0��3Sɛ��&ngJK�Ԁw,��8�V�?����*F�X�����-ڗ>��U%t������9�k
M��n��Ԣ���c�L�D�ˢz���ɷ�|\��6\�� �Ӵ�zMǵ��7
y������GJR]�hu"����#o��!ڮ"���Jr�`K�K�"v��[��>��2޻���]�z���"�kL4�}�L���=�?I6�$�d%���
O~\�*@�"jc}������*6`4�c�����T��nV�

z��L �l���=�1�]�oHw����ɴ�e^z�s�A�����O�Ղ��P����+?c�E����.�Τ�����xS{��+�d1�����VU���s����0N��ه��j I��|�:T�ῑ�]+^l�����A�Rc���pt1�I�2�
T�|�wG��ihl�T�`���%e	����߿���Z:Y�?׎��uo7��d4���(�#�Vw��U��J�ER���0|�'�� �D�Eܼ�*��#�:in%|�tz���}r��
,���Z\"�w���v|���i�9=�{Sx�:�`8���{��99iZ=��b�^�L�x�p�&�����O&m�^�p�2�S'���D�[��,]� r��{�Y�XՔ]]�@�0�_�h��L�q��x�!���)�K��h�zݙ��
�������g s�Tnx�X��ײE0��|����/������������݊�V����P�HHe0Cy��x�	!�yٜu/c�r���%��ok��v�������r��ߵ��;*�o�6��U�5y�J�xR5q4���훨����Q�f�p��4����u�0�G �5k�7�(��EC]��)K)�d_�n�kB�y�ɤW�����Q?!���E��шOg����D�\���ŷ2��t��h{��80;Ns;�%�uޟ�}@t���R1�a�˨��r�t�̨[�bw������ok��Ω��U��1�t%��������:|*�BgC����O��n�<���v�<�I
����i� �1Wj [	5�a���O4�*|c��~�b�~~�ls���~�E��k�?rTK�l�3c����h���Z �U"$�8�lh�0j#K���т�}�B�a_Ử�#�1�ʽ�t&]��c�=��f��@A�&ڳ�۠�kG�m�B\ă�7�]�Tζ-�V�t!��O��t��f��`#��j��t��׽���(	���	z%�w!�3�����*86�Zit��f#q�ڕ�`�ė�y*3�����c������E����L���e��ʠC6���n��g�Ќ�l�������*ԝ�u=ph춬�u-�<MX�E��%�@�:h]7��F�f5[�s����ʢZ���o:|���z�%w���n446x���p��$*Sa08��To��k��4� �N�34��墪s�g�Oq]nt��,\4�����޳�C~;/O�T9߶(,�f���̤.�?�̠����Ĭm0%$e���42������;����\	�1&����I�D�	���*�Q�ho֜��{�D�$�N~p۞��_}�ϟ�r�q�W���uLME[�4�W6y�n�nt������� .���FOoE@�}/�EϬD��XҕD�O��\���]���uѝ��* �������B�ۛ6��>l���^���߁ ��C���a��Ʈ��*`)'�n��(��zOOC:W��ȵ�@	s��#}R?B�����jphJ�[��ivDN)M�0;lsg#���TR���sI�Ñ��k�miut)~W���чs~���	�4<˼������������[=P����A��I���ŏ�x��Dr�( 8�^%�,�{�TS��*�f:�${\�&�G��pI�ǕA�^Rz�Ŗq'ͤ\S��Z1A�j�ϩչ7�4^&�د�6q��l#��
�����U��G�[�t���5vr%���X�ǽi� a�y)ۃ�-�����??�v�����k��r�tw����?۴QB�H<����p(��,�]��ۮ��xrQq���1Ǔ��d���".�r1��^O� ��C�|v�IQ�q��&�Rc�'����^b3��?
��c�N&ȫ���¤�8�h Ⱥ���nC+~�A��Y{�ͳ���GvtnZ��5O�<��3�U��u�N�+= �� �*l��{.�e�l~��o�_��1�
	�]�1wv>P��Q7�x���� �Ѳ��(��!�S�f���.b������aċ�v���G�q����G�Y�� B��V�������6�'l��B.���}y�f�<)3�(6�Y'�����7!�U0k�F�v����Zd_	�����>�*b�y�����#i(�<Z�kY}�v$�!�;��CS��z��P��2��4}y��C����
�ے��,F20��Շ�^�<޷��)OH���'�������=kd�#Q1�}<J֬�>']��V��
7��xò�v+�,?�,9��?9G����)��)ү����s�,t"ˣ�5��T��w���iڵ�M�&��b2p�/���1?�A�/�����������l ]q�_|��*��N�C@��A�Sp8C�)�6�nx���oʆ�\���V�,|G��s_�(�j9d�`�_��=���n⇝��D@��k�D�s�d��i�����ݶs<^�Gϐ��|1S��t)�O�Oǅ��0w#�׸�s��Qd���v������A����c�?{����EThN�chm��3h���_��\E�Ҋ���7bցN~��������Y����(�8Q>�`͉QK�@�hw�����	�ӝ�O�M�OQ����i#����"�r����,������_�L�e����L�FaVAf��ʛ���0�&�]���f�G�v6�c�jզ����	ў� ��{�T�g�����Y�Ky!_B������z�z��w����`�ǝ��ć����
͜����,J�'��ǳ38.6}-3)vWd�Y��Yb�6��Vd�!Z����Op�9l��������m��/��o&�_��S��#���]���d�w��+���� mܟ�r��ȼv�����RUN�6ۈ��8�'�
|1�i���߯ �><��&���(���6��N�9'E<� ���_[y����~E�+�$]��vC^��h�]��S��c�Nm��b��⦊���.
�L쎔�i_p.�O�G!d}�VG����'O76
�r�ǆ�#.�֒��ZİfWOlq���Y�@v�0d{�y�O@,����h%Se��;����bM�l#���n[���ζ�!7�ۥ�P�u{mp��4,��lI���.�K�u%OB������J�!e��kM��z�]���+7����&Q��y����B�璂|������ﶬ@V��4̷1�ܰ�K��IU��b<��C���
�k���=6+�o�j��<B88����F���Unt�9��G��Z���ћD����/kd˸D�n�Ҕ���x`�,/v]�e�;�A�A ;�pV���������l�Q���V�Z����}���p6�̪��G�i(���?+XtI#���Q��`h�8܉r���yL���/m�����y�5)n������a�����UeQ�z���[L��m)����7BΦ�ˍõ�;��kp��!yZm3G�)���Z�^�g<3K?�%̓db����n9	�2��L���1a����c%Sd���J�4eƅ�n1�ȥ�1	'�0�~O���������r��=0n��� $-7�ſ�9����|R#Q�['�0�ʔ_[��!K�x��r�,P���]C��ɭF�[3[&�w�I�N��ii�*I�F&����<�y��'�3 CO�s�]5���3��ZIa}��69+�1bq�OB�5�'V��/��(B�yu���s��mO9��n~}ދ�����󙙊��3x;���_[��1����M1��:[k�H����̯�lU����>K�e�ˊ�F����A��<.�ض}�H^p�W��v�X�H�3+=	���f��k�tC�;Aɔ����V�g��E<��V�˒#�j�3Z֢��x�RةQ�k�Q��S���W�=m��\�j���~=W̓zf���p鬭'e���O�~�O{�73`�s�;>1��1�*g��/7��b��^��M�<yN	�/<�����祺�?�B�~h�g��Q%�����Ns�o�o�Q�(�~�!���/ːR�[:	'�=�`�(�r8Ӱ�:�(��I�͜]�C�QF�I�UM-Ua�M>���OJ]i���u*���I�Tp�d=	t�(Ő����G�$u �D��G���|���QX}�x�_�+��!��y����\!�0®(w�0�#.�-2qg��'�����%E�Li[3�>��t$� ��|~'ՄR����;�QlK^�u[:��5�ѭ�����P��GjZɓ�f�";}v�|�m�Pgt����)x�Cq;��w%�,��8��Gw%�q��8�zh�w����o��[u��1����e���ˁG�T�Ϧ6�G����"�]�y*M���y$��`l"wl��bϽ�t�J����L���d8�ia�!#3���=�'�?w��Mv����'z6=ƒɋ^�B%IH�8o�n�8)T��e
0)�E�C!`�^^UN(�?u#Ȍ5�
�_�rD	D���oJ����#���F�
�e_��4��3j峸������&��Djx�=#��p� pB�,��	f�_!����QXef.z3(C	��eD$�˴@֊ �,ZN��~�	6a�zh����������I>  ĕ������*40��Vi����?���f3�9�+KAG���ߣ>�Q}�6��~C}v<�J���U�����w,��������[�+J�H�/��o�Y[���kd_Y�/~��-�|���~dx=���U��W1c#n{�%
K$jE��9h�t<2Y'�WP��{�ﯡ����#A�)m��Eݲ-�-p��)a�X���f��|��	�/e�[�߁G�rt��Һ���E��y�{J��}~U[rw��hc��x�7~.����?��M�V��=��pM�����0e���l'T�<CH'h������u7F�<�W<�x��a��dҽ�㨫����*����T�IgED�J	J�AB��WE�.]:H�n�B�Dj� B%� ߹xyޟ�����br�̙s��:s��1}�4q�����C,1_.'���M<c�D2���Oπ��<�hae�)u����v ��IzL������F�4�)���_t��ȕD�}[�k�6�B!�T��&��/��;lQ�v�뗽�t�h�sS�ɯB�'���O\��7��&���������j�s6-A�Uo���u�7]Ώ�[a_�sq�:��d�8������Tu��W�&'��uՃ�Y�����m:�tr��w�:^�j���B��J}w$|���/O�c�����4t��� A���Fg�æGݻ��/���A�Y�B:���	?��Wsh�,���|�O����`���H���sv�ɨ$�$L����Zn�N�����H4�z�,WN�z �)�Yd��vEA؏gUg��ˍ-H��x7��tfp��$��_;qz�^�)��wS�[�rT��V�W	8"G�!��WF�w�(�@~�}�	�)����ʳ���Z ?O_�t�a'���e����*��1�c�-���.���r��}q2N|�}y~�(��Wq�Ni��Z����$#"�߼�0x�ks�i��F�0���^�T��]
*&\J�����he} �qif���K냫�d��f�.�.}�+�*k4ig�d*�l������ �VW�����M��k�E`7�l���h���S�	m'z~QTGN����]n�:���1r��@�@;���$�����_&ku�/���;�Π�ѽ���+�t�$oַ�����iD���c	�y��[�}x\	����瀃;+������K�����tWf?4��-�ҽ�YK��3�jc�x�s4�yo:��}�=�[W����E��l ��j`�:��W�a(:p���Rnя<��iW�*M6yi���MmE�;�n@�\� �H�q��\8K��S�C8l��U۷�Ǡ�z��ӉP��h�l���5��^�Y(r��F����Te]����K�0�Y?)m���^��率���9�i�ژ��뒮c�F������
^��sR�[iXOWX�Q0�b�/ϼ�p��G�l�?�Y\b������ �X����_�&��m�%H�����>+��}�jn�~V�~��F�3���(���D�C3��lu��$2խMER0AJ^+�ё�8o��U1t �`ݮa��:�穽�v�N�i�|e��閘���~�� �>�Ǌ���>�TK�T�����օ�t���s,Wi�.�ʯ�$�q0��o�����\W�n���1�?i�b����fg�Eq�!�����`��Ս�+\�::-δ�q���O��#k���v;�]t0�k�?������(l�0�O^����m��.�n���2864/�r�����TO�WM��Ik�w(���ۍ��[Zy�._���f��¡4�J��-��&�	��Y��������}��-a��{��,�T�`�ʶ�I?{��C�o�٫BNv_V���;A�}=l�%:w�`y3ñ��ŃJ��:���`g7���&���]gu����
v�>�+���F�j�<L�=�N�笛�lI��W�Rc�Е܃A�Zm��5B��v0��G��j� 8sY�x;t�%�������d��N@��.[���,0Q� �*�/�!��~���4��q��6úI��g�K��P�V���j/h���s=���^E�'���Z�GGc��gǬ)�/�F x|��_��馫�O��Ё�Og�o^�|�H�)+������2[1��D�i�;�0��J�*z���'���a,��	�{���0�m	c�[W���ͳ/𕚤�ؤ,-��cb8Ulg�Zk=}�%��,�N�n�����f	��Jo���\�ġ�@���0#�o}��/	^6��O
 r̚��V܂����#$�����ט�`�K�Jǎו^\��Y�rB��C�D��r�c��'���m�"�8�O�U�=��~ �#z���僸�o��@���8�;��d��&�^Ԋ�����=�᫝ʰ��G��v2k�[�9�� y����i�FBģf���(�����z}]��;r�X1阂ם�i�׀�!�*㈲���|�q�4"y�, l�����*����]LX�\~���m���N���_\����r@��p�}����`�HMǣ��M�J�*b�_��=F�+�%�Ux}��B��A �>JfGػ6ALJ�V��~��Ά�t��7TgGt͏�,�s�1)*]�\6��쫙 ̭���t��#�������A]Q4�8�W�Z[[u�k��ir��F�.�ww�$�;��a��e���l��w*�4�O��Rޕ���0-lQU��*?#�p����&��s�/5�^b��z�*3�K��w����
��T`�[��nV/ܧ�A� v�h��&��nv�U��Ȼ:�Up,`����k��
�Ba_]h=*�)���.~݀d��M�.�&|���Uu�\�����l���PX�����脌\���o��O�H��X\�Y���H<NCII	��y�^��5 8̚�����C�a7 ���u7�!���!7�zt���7�>�nf �y�+W#�3��rƭ�W/f's������'�åk�����uwC�p�~������)� 1���h�H�:�`�� �n�I"2�2~3������.#��I�����F�}�uٝ�q0�e����^<������g�3�4]��楤܄�v=~�a����d:L�c���$�R�%�;]G�p(!#�˥�pd31f�}�V��sY'�������L|X�j�z���ex��	�5-��&552}�m�tө@¼��6,�2q�M��b�~@�i�P�-;~�ڿx4�_F �M�������ć'��2,��f��=����O��[�׿�>x-CT7�������i2z�_8�z	�}%bB2Ew�7�y���/�B�����t@O���_�~7����/�k2�d=��=�dG�1�(@V6��T�f�B*an#��z9�/ߥ���K�v���l�G�\�"1��U�5*8.�3��r]��'��K:�W��Ƥ�>����S
�X4l�h�1�����1A;�g�\��<��7���߭ߍ����*�8��mᓓ���0y�\��*��ۛ�T+>(��(��Dy���,��o�%���/�U��]�p�x���L�G �x[������3"|�)"O�_�+�K{���8{�-�!)�"nk�����f*� h�f����@b��!mrL�srs�ʇ2���^��0�叽fݢ�4�)u��e���g"R�-f�~٫��/�X͔�|t��.�@��+j�#çt���l��wbw���l��]�56��2%��Zy��6��m+X�!�.8ő	 � ����T"3�U ����v�h���,D������3QQv���n`�{�v�Z�0�%�t���R���W9V.�V+x�Sz��h�nrҰhgsuvu2nX$�K[�c9,��左�Ʊ��u�ܟ�VR.�H���S���-f�'�.��-r!er�l��	���y��0��;��0���Μ��I�!7�̔�z�D�A77F�i
ރ�'��	�3��N���2�i�8�� �*Rw�������u���?���v��;�9�,��n<���3�#��}����M��������j5�����A9��=��C镕2j=&(����e�'O�퍔kv�P�[�w�JF�ok�yH^P*�땭�U˽��l�Y��V�TA���FJ�� �^���r�l��T��lݮnm�_Z�h��=��I=҄[F�� `��w}��t�J+@2#�~ -41�--
�X�U�T��=Y�Lqv6�ߧ�Ta��5B\�ș�����2���wGW�p�b����k6g�����]���q(B�Z@@@Tn��t�{ڠ�������]VTƴ^�7*��+6Rnkl/Hn����©]i�~Tn�=zר\���-�Q����+��Anm��!F:Z%��a��u�u]�y��jS��s���ع���>t7~��YZh�"��~�����ׂy�PƺI��(��|����S��Km^ړO-LML��X~!䀽�����cG^x�x~�I����b�6w}q��P�k��k��Ǐp�����|�W����p�P���A^ݼ�`����L�u�?�;������j�l_�җIN�oO�$|c����I4�8��SUHr�'��l�$��y��v�v��5�K+*��ߋ�PG��,�cW��_x��~�-�2¢�b([Օ�5�F�̸���W�a��sǋ�h����>hr,�U��=BO��oW`���S��<]���#��5�㘤��_��t�l =��,��}��GMb��^�_B�*(��j=�����jW`��l�;	]:t�s�V;&�J�Z@��}'�|E�T:������6��BH�|�h��H���s?cOz�i��1��N��!��R,? u�j@�w��uQ.�������yZ�Nۀٌ6�CF	����wc�nI�jvC�RK-�ε��w��Μ��9�̗�o���L5���|��<�4S��Wu�5�`e��
��VIl	������nܙ��cٴ����L�]��R F}�40�Rs���O�B~}1'ے*j���ZJ�=["W�Y����q�6n����v@u���s�����X ��ia�6�a��sNsC�}s��}������"l��=�	ٚ}���/�N�M�*���WӅ|��U�!��O^V��fp�&esR�������F�2����=,wLȯ���<�8mAI��H��B��V���w;0Dyg����D�ƣb����B�mo�pr&v�����q��
 zSb�A�5ͫ;<���z�5ވ�6�=x�?���[i����;v��Ы�S��(nA�o��: 7���I@�Mm��\����,����U���SG�Y)-�m[C��`��D���K�~0�4��^U�?���5����ra嚻�Q-�
�4��U*�����7��wxr䵝�+e���%1y�!�V\O����Q;��>v�baS}%ı,M`��c�ce��n|���o�K�fI��9+��|.�c��v�����M+G���d�Q���1����QMt���Px
���o��ǏM�q����	�����*/�R�J�M�x��@6�۰�%��Gq���3�'�YVM;5��LM��s��{.%�◫���m����7��ݎG;|��?����2v��������/ΛGZH>���K�3#ڪ��~lJjJ,��o�������M�p1�Ƿg��3��C�	N�Ya�jjj�%/�.��~l��b�7�����^iM����w������i�Q8=�� Μ0$^`��Z(��X��CIJH̛��ӓ�q���Č�dQ�)Uق������5�=��-i���KL T;�ʜR�;���>�V���1'i-?��9ױ���-�]�����f[48]�m��JI�KRF&a^k;@�«���3<%����Ro�����t�X\�{��i�A>1�O��>Й<�1�Lm�w{ǭ��-tAb\3ڄ�0��:�~��b�GI�j�d���+Ű��":���r$�&g�&���3����}_���c_�<������2�C^4Rhd��0Z�rH�YYΩW�d�6l�v�����k�}���V����[�W���݌d=wn*9lll�K����C�@7�,��PG �g����PKtu�ʞV�Yl!7MdD
(u"ѳ�I�M���YgX���H�L��I2������R����A�i����$�D�����O����=<u���rw��b��r�ތ�z�2b*	�	{	,p�|�WGKYU�����nŭ4�<Gk��j^�W��ѷ=,K�Okj�9�>!�7.Q�CZ��,&fI�)>5;�w��B&JT&g "�����8#m�ӥ90��߷z�����vR?�?��l�d��K̳H\2Z�j�튖p?��9�\�9�;#P�NK����D
b�(�v(t���O�GVo�^V1W\���l@Pv^�c*O�Y{H�����U��H��#+����&�v��?��{z"rz0�g�08_K�ʻ^ĳ�� u��z{���ߠ�$�
�Y[�Y��5T�*�}��5g:��1���{�т�ETy��m��X�$O,�آ%
*B������z��+�{=X�޸�5�@�#�]��9����1M֪��᠛}GϤf�_n���nOʳ|��Iq�-��Fջ��k��<�J�7q�
)�2_t^k�Q�u�L>��Qs7��c\N�0,;���궢�#!���#(I�p[o��Y()��Y����@�Ы.�x��{T�;�F�8��W��旡���H�J�b	�5�����V����沁)6�2W������Ħ]�e5R�K�����^�n	KHH zBtM|�%���פF��T�Y���E���%�B�0�����n�27b
�����D�!0I�h�O�[u,�ٻi��"��xc�ccxPni��t�Y:o���f��Uo��5�缵>��g?͡�\�8`�>Ojx1���>H�a6�[�e4��g�P3�0��JC�T&̆������n�qv���j[`�g�y6�|r�P�tn�v���c�o���F��mmm�-������<1�EV�D�q֑���D薾0�.6��w�	���9ۭ�`��;�nM���qF?=�g>��h�j�1�Y����yEb;��l�n�xתeE?�LtB�a�2�o�����<Gq)S��b�y�6�Ƹ�ZO�b�Ȩ_�ـ��SeQ�dM������kݏM��t�Y��L%Qk��M�?�8~B����x���M��}�._�������k=(��tmAtW�<������^�[��CԔm��ޞd�����p8�A~gɇ�Hj1���Xzmv���~9�<� ������*F�d�96�8&�ב�TΝ4J/�*/�7�>�E�V�U���m�Pߙ �U�TT��H��dG�F�m؂�h���짼��Uvf�^{[_��t��Z�7_-���O��������
�:����P�l%�J�����0�ø9]���dsP�p:p��� B[��sI�k��Q��ND�.����|\v�S<�p��� � �$3BC�aa�"O�dUеh��:Q�J��˞9�-��,�$B9��`c�a0z�;MU���j�jr�+��of��z/T�g���������'��j�8�2ǡX��������\��H��|%^v�)�����M��՟iF��f��C,���Ӥ�xd%W����D�(&9��_��qt��Y���#�n��R1��){v���g��g�%��<�;�ځ���%�[���LO�F�u����}�� ��I}L>�K��9�Y�0}&�>ǂ�p;��|��:;xHu[����e@9���{�,D0���
܈l*i��m��i�HGI���r8�6 �X�c���h%iQ�"U=q|&1z�ˑ*a�2�#��k#IP����*$Ȗ;+�K�pn�����X��$��T4��� W�����|@���H�=�"y 'ǥۅDs�>E�D��f�f� ��2����OU,d��* �	}4!9;^rh˾�v�0K��sń�2�)A����\�qn�:�dYru�n�����c����C�Y�'''�P1�<�����*Ae��^��:��^���IJ&	�M���w$\�&�%T�Z��^��K#V��oN�p��,�޾b��+�Br���5����1re���F.a�Rp��ׯ�'���}����.�c-�4ຘ�j�IbWӳjt[�J�0�;��T1Z�<���i�c�3���B#��%��g��6���b�61�D�]~Sk�����2T�c�<�������d��=��"4��Wi��R	؞X�<a�~�)l2�r�r���̝����»(�JR/���t�N&��3aD>t�`���}�*M�*L'���,4�"�y	~T�%Ҁ4��g��N���U��ER[[r��Ź�"��xi�F'H#ևܭ�k�}H���%�'�'�j}�L�G����.������Ġچ���\�o��b3x�X6z� Qߑ+if�~���sR���%:�[�+���M�g�JmZ��������3����h���pg��j�v~�r��'D�32�%���gڪ}��hI�����At�n�֤��eu�������f��sZ�:|Q�4�@��:{xH$3U�~�_�O&�15�����՜m���WϏ��;�����;��K��;�s�A����^�7��7����&T%
�j�7�6�%J�"e���l4�>W�\ (��a�!����nL?�U��/L%������e>��>Q&�{� �����j��lLgn\��E��*W�{6!�����Q]���\�P<;�F��ʫ���-����		�r�)�w�z������v޷���egr���928���Bvt�7�,l�����N��Α H�� 㪮����c(:�'�y�"L�xΐ��p��YU0�rdy>QhCE��c0��^t"���sۑ��)�tT�L�m�+qf�j�_f�G���v��_���u�z�D��I~H>�2����?Ҩ5`�N/����8�&����"g�;K��.!�kM�T�4Gls��u����B�l��T��lu5\���_��:m�d�"_S���>�qM�cKs�Q��۱�X|����J3��8�^Y����L��l$Q�`��؛?�R./;��������+r�y0~� �3�:Z�MK���e�>?|�p T�4��;U�WI���n��n'IH
U�����o���@ê�]NL?B�~�(Jd��s��_H�#�|=�B�%�v�Uk���?	'^Ř/�+����c�}�5���S��˟7dy�Xz�[���L<��1��GZ�>�%
�O����xK���/�;��2��{yRӲ�3��2�X�����x^nN"Ԭ3\�yˉ>��Xb�7%0��D��M��6���]i��V"z5T^znZ���^��k�I�┌�#�)�n��/p��m�>ݝ�6>$��iQ�~/�'��)�;��&�ؚ�qi���������Q��lZ��em���(�7����(��B=��zz윤����~	�r���n)����!m�1 �������$�wRs��R
��Z��J"W�&�g��� =���*KX񃒉�Dm�U�o�y�R�3����m5�zv����޳�4�4�U$}�=Z!��!T���N�$�7r��B,�Sv&J�J��́��ܩ~�uԽɉ��3���Lq9џ8|g0�9�3��9�_Bp��!��h�(�_��.�U�<� H�r#�̞0����Pl�Xt	�
��#� �Z(H������ezO۹@ �E�������/�=�F�w����d����=�3訛������,vR��i�~ߙ��CN1+J�oO �뻤]nX���@�n�q�AZ%PY����A�-:�v�{ڊ�x{�C�M!L��.i�
Kž6fä�
�o&�i�Ƨ��s�Y�`�p�\~�1�Y��iV�2��M�����!�"����hUM[��q���%�͇<�Q�.i�v��1]Q��!7*�����=�m���e��~Nq�����!cyL��*�e��p�DT���}�v�Dz�u4��Z�J��m�K�J�L>o/�	�V� ��1D[�t4��f�ϥ㻾ejm�+~��뗏B
�O��a�+J�<1[�i{��\d�揦����@�:�5܄ML������~@H�k� qpF�(
��i6t�w{7����C�M�1)��C�1�ZA�ҥ���i$Y	�e$����` ��3λ������F~v�E hb��B�8W&*8����ɛ|v�T��](99rR�n\zZf��*�2-������ĖIX]]��.x'9K5i0�i�2��DJ�D.m*��/Q0de���¯���`}��}v]X�Ў��'��Ǣ���͈�p��H�h�>]ZZ���Vjx��[�]�S��iI;q�hgυ"��O�~��_�
Z�z|��S��[�UhC���8OI9VD̸I�����_�]V*
D��Q �]<�p�����I����7P�o�#.Ck�@|� ����֖�9J�� �
.G���n��3��q��m�ȋ]�Qk�d�A5����~_�S;�h�_�'G�y�J�)���N�?��Bn&�K�}`�be)U�Bư�@�V&���[f�ʌ�p1��C�ǁ3%^s����PN�{��*�Xxi�j'��!�.��b7{��G��*ہf<�v4��`P����D��7���sϳǾf��v?��M�.K$:��5��,jbFn(J)�BR�J�&O<!ї۸�3t-�-dpQ� �ek!�`hf"j8=Չ�aQ׳�f��9����o�&�y��Y���&r7X���K6�ި�L6�;@���&	������eq �4��+�d(������=�j��9�u�%�r�}z쳆`K;���?�unv�k��t�s�kS�fu%jm	$�_�7��9��վ��JBpr[��.%�g@4�z���x���s��]���n�]������r���tc�12m��Y�M���74��툪7rq�A�慨@�)�mЂ@�k�� %
x%�����$�=l�R�-5��аˑ�Exࢷ'��^�	H1�5�rXڲhWwB�erҍX�a���nk���G�v[�(�"ۂ�fP��7��*�1R�~��1H��	�/��p�jB��� .�\o�z7��>&����GW�;��h���y�Ѿ��=Gk�����P/3s\����2 ��5�T�`'}����{�@��1~jƾ��0�*4?}��Q�u�\"d&X��;��{�C�N��,��a����4b��d��u���A�h �ZR��x�ڧ�<3LX0�L�`�{�D��� ��E~*M�G�4<�
ĵ) =6�T��ȹL]���z����v>��K���'�#��'�n���>��]ZU�K�Z�v��������ِ*�_�[1�t!�J� �W�r"�<�� �BYi�c
���� ��_Ly$�A�\���n�l���e�Ӫn���5Y0N�Ά�y��D;�Zk�C��`��p�Qe����	%e�0ݜ&�7��}>��վtJ_�mޜ5Zm�8�[s�����R�k��]����a��d�A���`�r[���W�\�P���k�K>6,.����h9KX������A���AG��lm��`��e%&�+�N�����M�_��k��= �	>���/��R�ݵkoM^;q�j�R�%� �A>�)��ùL}ِ�u`�Ì`zW�.�6LuxcP�O~�i��!����~gO�2�J_����_���}K=1�\FL�l��5q�p�bd�o����>;�n�~!��{�OM+����%@�^-Uh���OOl��VݏJm� � �)2�Fz��r�i��Z��@�2K��hW�#�I��׈(q&63�gg@��Ci8T�t�]_��"8ug l�"�W�	xD�f:Ż���3}����~���b鳪�$���8�f"�2N��	����g���þ�ЍA�P��]��i _- _���Y<��$ew�YŝWo���L���TG�ϖucD���d���1Q3�v�B��C��[�ò']��=K���2�r��0�ɐ��SjyL䄆(wWnGL��1u�� 1r�9�I%��3l�	{@)����A�ԎQ�/5��J�0��Y��#�!��p�Q���Hj���P��%i��#��v�y�v[��2dX�����1�S�%�T��7��ӏ�" [�nH���ڥ���^�pt,c�c�_,�`��Z�0�߳}y��`�;1w��������`K� �@�c��]9$J����7�`F���Wn�~m�"kl-���©�#hnY��#/�4�Ux�%��]S(���c -Or쬊��j��fE$��w�wŗY���A�&+>�,Rf�E�K�!���P�]�ҳ/xM�>'�F^�{�~�k��9uOɞ>�d]I4I؎o��x��9�V��ܮ�hS?|wd@�j�̶�k G}qB�8�Uj���L�q���#u�v�{\����C�˓�4P���ż����B�c����ӛ�x]h~.�`���J��2ွ��9$7�L�IL5��G��\�o���P��gj������z����l�c323�o�>����Jʒ\����˃��,��u��^�XN�W�K����?����h]S���x�Db(-K�ޡ�]<�=6�
�R�;52�ӚPB5�x��M�v�F�=�	�[I5(|��~o4��ȝ�Y�ԏ��.Yj��ww$��Y�?�>Z��Abqdgȑ+7o�z�r�ʩ�S�e�䆏Ys� �M�K&��ʇ唦Ծ�Lhn!ќ�y����~�5$	��a�Զ�x&//�e����ߗ�w�=e�K�f� ��S��1AMh�fPs`����f��~u�����,�>/ e`�U��5��S�3Fa\��wgg/���]���Dul�{~�X?�Ez�w�^����[E0�V����y8� �&X��DJ4�_1KF�ti==J� M{�յg�"�R^�V U���$lE��6�L
�>c~���H85=h1��[�'��*�v���t���n�z��)1 ) `R-��ٕ��^����Ԑ��Jנ��:hu}�_^�f1�BI91�m�x�0 CO���>U��^(��3lԽ��=����{ȄNCeee��l-�Ђ�;�b6X��J�O;[O��h�ĭ�<X^.S�'����&���E6p��ԑ.#�3&�s	��Op�g>-���~��a�("�;���9��Ώ/M��i{{o�����a;��ڑ�F��_���x�N�Ўd�e��U:��8�E�)��8������%����9���>D��L�є�&'>�ݰ�8�M�X���?��)���>��*.f���E�j�!�BU�۟��B�s1yh8��ں� ��i�y�~SR~z���lR�`���ZLڝ�/�����#- ���1���c�N�-�&nL��dк����\�>R5�g9<����Nd�]�:���	R���rMu�H�4,�s������q2^��#I�i�~�}�gM0�#������+��+����$ƍ���줌���$���$l$���i!@���#�� = 6��Q:r������^I��l�{��r�G���J�Ԥ5����[|�q���m�2���	���B�a�%�ZX(Q��٦�ZPe)��E�!��r3_�i9%U�Zj6�/)od3���`pw���X�^pl�	��]��Y�5#�6�E����S<w��w��I[��[�V���S72
�����ho�=�� ϗ3�:�>�\s��b󦰔T~�_Ϡ5$�"8�+�X�~���|�E�?����������~2^���3z��N�6�Ա��O��u��)����}Z�P�>��la�p��Z�m�_�֟b�e�h���i/���+���=�ӥ �ձb:#�,���j�{zM�<�������}��x.����������N�6����rˡ�Ko᭵�
�OlS���NF�Ğ�[���g'����w�����[VWW����T�P�ؼ�|���2C��93��b����j�)��//���_�K:_NMM�qtDC���\��_<����<�Vbr��X���1��y9�/9E�-.:%�u6���Pմ%b���ǖ�W�dWu���9M����*o1�U��x��2�fFʩ���5F�Ц�A��e�8!�;RiʯE��{�D� p>���Ǐ�~�r�$R���	�i��`���xt���ϗ1&o�~-t��z��I4�}6D~ǃ�¿��!�Q�2��3gơf�"�n_������x��:��%�� ͈s�j�&���Y�?/�'Y�S�b(���+p�o��bdG��J���]��,r�(>"��W�[|<Ж$��Bq�c�'�r��o�����6R�<)�V���DT����P�[z�`1�$~2���	,ԸE�W8MX��ʊ�@ٮ�<;D,��]#�`�������vh�yx��ٹ�i�{����}�:ٜ��!�C�6�
.��������x�w���#��j���!�nZ_��YS�{}_��Q0Ǧ�r��sz5�ݤr���u�}mv5�5,'�Wrsrr���������oZ&�d������]?ʺ�|���+!�T,���:��{i�s��暍:�=X�`)�Ơq����|�N%5Q��=[�3��[��1L� �);�V���_�
VI��[Db�-o��5hK�nN�ᄁ�������J�?��.l�&_�c���V�c|���^n��W+��S��|z�S�����O�Є?c�����7qD������y��ښ�c��K������A쟘c�Ρ	8e�lu�W'�*���P��B��FȢI���#��g�D���sFf ���l�v|�9O��6���W�!�����Ib���9&۶����-͏ݶ;��K|yy9vn��3�rC��{526>�׿�"F�RCz&����D�{�*�;y2�u���$˓�/���IzW���P6i��9�}WR$+�{�YZ	W�XZa��M��ua�w��ӱ�/~-t��kmU_#�~�ɨ��D��������:a?2�f���\�k��wM�ϐ�l�;%���6!���4T$XLRo_aE<�G�"ot�/_�E�Z�aº A9������2Qr?�������L����+�w�ݨ��_l��L��ƯV�Eb��}=8�x�=\����Ɩ�����? R��{��PNX|n��z_�	ԶV�t���3���}C�b8t�ѭ'�Sy��4�CD�o?��#���-�Ժ*�u��ω������=�^yJfF�X/g��s����3������@9\~Z'�����l�s�(;���g�r����n`u��]�=Z��gBR�v��">��;�ŋTA���l��9!v�0���������7����:㊀��+�@�J,C���o��e�c@Q#��������
���CX�tss{�Ƹ/t�@7��L��4�Ғ	moo
���6���
1����Dg��eA�_A�����M2��Aj�������j��&��}���`����6�&���)t�ٙ��N]�W��_u�x�S���N��ǹ�Mb��_���=5�.�����'롽� ��ȉ0(�����q���=�mT��l��`f�J�����������7�7��M-Sk)�a��O��&���L��(ݳc�I�܂G�����t��7(}�΍�3E�Q��V'�C��Vg��?�x�����߳�`>m`�������|�՝xƄ;��w����.�*��/}s:1�&�J[��C'���U&�-�|j����$���-4��.�&1j��$T��"~�Z���� h���ׯ��d��A�0��������à��\g��.`��J����x��s�j�c��v4swr���ޛ�:t���5�#Ф=������ç/�@�����m;-����ĝ���k��'55�������-����5�;_g�?�K����x�l��E�MGG��򣽯�
=A�D�|kLY�UR+���+���P|�W��v����m���,�@����s/r����KK�ߌ'�BB^���W��-$��Y��K�|���:��g��mq�/����;a�J�c0��7U 7bqm>i�z��V��m���Ǯw����Y����A%ї�0~��k��7W�L�X�����O��9wmVY~�tO�^jﶣ ����/���DT��� ��D��Ɍ��#��D��Ћ��u�Y:34Zl�A�r���M�IЇ5u�;ߡ\����C�l�������Dog���_/#PәI��,O�\�u'$�Ͳצ����\�4\b|��'3�.l�m����w8�]pCT	N��:��KKK�L�G�~��&bkg�&�3�*٦`��O���,|_e�5'g5W�E�z�U��v�%�x]��}P�K�_��.���@��zz&Eµ������dÉ���6��Z�^r��%op�6R(��|lx�LF�0��� ~�DO˹j2A��}_T�!�6S�1~@�/E21��zK.h�G���Q�|�c��@M �m�Y%�}��db��������3)�?�31�0!5�]�l�����?��ά�HWCD=�����x�����w��U��Id#]]�	~E�xori"\k��P_�+���`6ր� Iכֿ%I�,`f%++�|� /��{��	�,�)��\^^^�>CF����Yl�`�>��u5G�Y٪i���T��Y���+l`���'h6@����9���]���R��Ĺg����M��K_�C��?;=�Z�l��SK^{-��zŷ��Z8�bVʌ�~-�E�K�@\k����V##�y6������eα��Xz�$i�����h�]J9|�k5Z���=�}N�}��J���b�I���O�س�9�s�عf��3U����;5�kB'�6F���G|��A�6����-%&���A�8Yq��3�m�����X�ǻ{J�(��o1>�"�q����*�	��F�0�	d�����=~ iA�������n��l^QH{�T_6�����m����� �:߀l
����=ON^��4�<8������g��&�HRϙ�!��0�#/D��zoL}x���0�����`�����o�>�z��{�	�@g�]`�A5V`@����|f iu=�l
�R�
w]�������fw�@q^K��;e����ډʴ禪�N�8*�!�c8r��`�%��o,Z�pR������YqQ�Q���8�[�%��Z�3X�w�����2�����|m��%j���	m"S���o�� ��O��h)>&ÈY������к��f�/�:��F>�8
2����ӯ���,~1R��r�[�i�z�ީ�����RGs
�?�>�砼-��mA��:�/���Lp3�7��1��Cj1	�^���k� e�:66�����:�
�s�#~��`8��ܬ	�ZzA��������ռ��#~��Ǎ����	�>�9[ gyo��|�]�OS	wf{vq��օILR�,��ٽ*�z�T0^����>�c�~F�(|��އ(��	cu��\B����g ��r��l�^�v�)�\���б:#�-�դɍ~lux��<�&ծ��2+?��
LPI������o����+-{/�]���3p�Ԑ�Sb6>RFd��D�]Me��/Іn�����b{__�,��zVxP��j��c�ɞt<2�J�����u1V��r7�mbO���y�;�{�u(�j�w� Ғ�A���!P�	:?�E�F{���?����9(v������,o��Ю��dA�S1���o������rR�&Ɂo|4���c��Ӽ��Ҩ6vV+�k�H���
Y�.���"s��8	���@�[�B�g�
���{ �C��x�,�F�݋g��wQ=_����ZK)��D.���Q��� �@���)/��:h�@x��]ڮ��Af��-�^��؋�m��4��c�f>����.���l�!_���c�����F�������
L����l���W'u�2#���3^����Ϸ��_�5<�X�m���5v��w�3���".�Q�͡�I#����Ng��`/Pv�p&�����+�a�Q�sy/}N�i��������1R~��S�6���J~/r�VF�3Pô9
l�/K��8���j�b/R*��Z����BK���S�lu�v����]T7�2(-�{�0��J��g�9�ˑ.�A�������H��Zp��J�p)l��GL@�e�>��P�{���u4�8��B�ޛKX<l�'�u�������{�yAMT�ݺz��M���۳)E��#;�Y�x�u�z;���x���T�O3�zG���o���z2WP^��C�	��=�q���>�։��ڒ%�'��t��68 �u��e��rj��ݾה�
�Tʣ�6@���w����dojY������"�+����D����|�.u˫	K!�l�=�8�=�*9�����dT�9���Ç���l��AOG��m�W���i4�)i��S�W"�T�]M���������۬y�V��.��(�S]"��[(��8��޻���B��2��$I��BZ�Z+���JTō�����fi�T��I8��H���?I���P��Ɠ���c�-��Z��a�(�@DB�CZi�nPRZrhT��n�$��A%F�`e�a�n��������%�x�l�X�^������31BJ$���ƽ��Hg��������I[�7%�掸�`�_8��Ғ�#�� �r��4�	�b;�~x8(7)����Z��V�O��:�_s��!11W�>�Uu��l�c��t��;��*ãS<�Ӛ���5�'4��^�ϾS���'�f}��R
ibg��s���	vR�����L� 	�[!;��J��I
�Vήf��I�S_�ǝ�D�vUf���	��h�����j��u������h��6h���e���D��r�F[�C���5nv����J�%���)�p�(�2�8"��/M[?>�"Sd*q?_b{�,T�ض������ez�(H�>?��Y6��]�����r���O8?�� ���Kxjr�bǓ'߂�an�U����,����gv�4���q�~[R��R��q�����9wt n�܏�q����Z�6�֒��y�>�~ڸ����R�;+�{ �F�x�P�J�>2ho:[�2���f��ô�:��2c�E�F*	83�l{3��M���ن1&�u�7�WQ��E	Ѻ19� �v�׈F��%���'�[D��sz�ģN' |�ǛZt8:c��c�v���`�N?�;ڽvҢj�S����E�=���g= u�Je�8�Ѡ�&�Q�-�E��&�ə�o�{��;��QY�����������W��X��=׈#�X�L#F��L���0E:��������.���M�4���']ϩ��.or0<������(�!�c�-�m?���C�nh�{�6p	�y�?��Ъt��g������4�ӇL��O���ޙm����^,��zt�joNu[U�a1$��{+�uz�	)5�N{��(����M�<�ڐ���{�ȇLy� q��z��׿����UD�X�{L�"��JA��v%7�G��]��gk*�DM�Q��="%d
~���s��9�ۘ�e�п�����f`���O =$%##S��61�v�}�Ȇ�� � ����KQ�eq1bfo���v�}�~��4?[GvEF�~��`~n2B�9���`�8Uؓ�7�uDb��z�i ��	�KU_7-����\U����Y�|�y ڋdfa�ilBrqW9-t�6����qm]ݢХYc�L�}ι8R��@�`����a������|> 	*}�t����;.Bs;���c`t�ifؼq)�fv���(
���}bbuky�L,��)u��b�Pr9�Z��[��rN��iWTD^�A&ehhX�cf�4���̼�3���6�Z;vȸ<�N��Z���w���j���yh����V�O��P�r��)�)λ�)ej�^��Y{��$��S�z٭4�J�O���Ylqvm�m��� % 1Z�>���aIU!���U��8�L&����->�f�(�����ZV~�z���hl�]����n%��V�<p]Hl��W��o4xeh��P��{Tફn"���P�� ��g�g�j�K��-���3:�Z'P���[:�6y���T�2���[�D"����Y��e��T�yWtu1>��TB�H�Z3��x�"O��� Gy�:aZR�?8�
�ѫ��7��y ��Y!&��������>GGJ��陑E��	c�6��}	Q��C{��=ʢ A�@QeUK��t���9^�2A%O:����`��FL����/�	Z�h�͝�یfES'���rt ��G9��Xc��) .&�ieo_ ����n�b�'��9�~����sw8,~����O����@N�tG����x���Լ��\�cߓ��i����r�����e�|�h���5�&����?�F���<�Ydu�-bS�ڬR�yU�E�η�!��PY��^F���}s�~1�op:U���f-�c��Q�!�qYa/����(eb��_u0O��L_D}1��T2�ݑV@�-�MDI<�0d~���M�"?�Y
@��X�eȠb��C��a�H���I��;�>�bAL��d	_U�����k^�4h��ǁ��n���f~$��{�I��7լ8�ޚ�z�:����P�~E�=���[J�~�vb6P��dԘ���Ϙ̵�r:7���}`�흾F�(�_��8A�cp�QU�����[������U��-�j���!��0��m��$��<q�`���Y }��cP��sw���:y����1�i��nM60�'�+pA���@X��e5&^���[���(B��ZG�yQ��'�x�rRטXe������i�ǯ�r����ȁ�4w�g=��p=j��a8JC~d�kk�b���"���&��pj�%�r����;��1?֓��z�t�A�ᾊ�L]o:L&����K�1��22���"K�x$���� ��Xf����d�	����>.�|���39K�%>+W�&�����sG�9��]����b(Z��C�]�F��(R�C/�U_�W�wˤ�I�3}n�l��t~f���S��\[pCĥ�g���{2��:���Q�Q]2I"/gba����Δо���P}�qC2j���I�HE�e���_�ϳ'7Ż��͠��T�b@3jz�'_"��୮ep;3U@� ��;��o�+�l�]�sI2E�o��1-:�-Y�F�<����x��z�w���Y�����+�_-���0�$�2H�����SE���mk[\��k�Gշf�9�yл5u���' f����b�k�u��^ . �1�ǭ�t��}�Խ1��A���b����Z������x��aYCS��ȟ��IV�/�ml���K����+{��~�]���ѕ���%!�y>4~�T}�\���kZD�,�d������I UX��*a^�q8��}d$)����8e|�c�VYBO�g� �v�|'��t��s H\^�ZT0�G�FJ���gK��l���:��'�I�q��>����95���Z�4>�Lm��(U>�q��X����~8�rq�ā�q�ԉq��jE��bӠ�¿�}�Şd.����x�v��r�������DR����N_eϜ�b�������j/VVM_�X�X~�������8#�F�1}�楩��M�	��B�Yu�ɯ��@�ڢ�r�����s��6Ͷ_&��AV�Vվ�O�ݴ�k`�٤���)��X��A+��0z�Q�0P��^H1H.;�Ś�"����p�oT������2�,�%���3�p�			uI^�|sx����ŕ݌X��7��'��F��� *q��e/ʟu��$�)))�VK*h���Q�?��P���=|E �kf���[GK����&�oR��î�9⹶�|m7*�a; �J�9��n�z��"�3�/c!5�0-�j�c�®1���U�'{�P_|(5{��x�����r|�Q�[��H}R�A�jj���У�Y؋ч�ɴ�����J_E����+�Ȫ{�v�+@9���2@����^\��e�7_U�u�S�f��Alg�����G]Ǥ�4E�������3�{o��M����-���/%E�wVd5jGzƚ�9��~8,f n�*Z�/�`@�<ذ����	��N~{z��(z�}�<��$�z��>��%u���G���D�ywBi��#˳h�ޑ7�*�ɢ���T�%1�4�ш�׷_W�1�E�lQji#F����?M�R�S�ǡsr~<80p[��Usdl��5��	�7o΁�=V����U�®��8@
|���pK�%&�;�cR��j���w��ܷpʪWG��9�/�R�I�]�w��\4) `ғ).��:LTуY;�F���ր��Y�r%�N	7ܑ��D����<٥�P�i�J����R�Nzw��.�1�ҍ��ߜ�=�j���0�����Ӎ��z��7ڞU!��3Ծ�%�4��I���V1��N�SSt�bdL�F�s�װ�
�7@V�l`4���H77p|~���inV��r��jaYY�P�vE:R\p�����7�2�_�jip�U9�@�Q�� ���yʗs��=<1MN�#���e���<���_W}�ǘ��z���K��&�^"��
��;�Bd����JL��$
9M���὆g��p�n����l �)���t�� u����~�#���Y�E��'�%�PMs�S�u���$"b��tB��::�Vۘ��y��Wu��*sU�;��_Q�ٳU8�S���_�3?�:�LQ�w���f��[-�e����p�ˢ?�zs�?�	��kz<�vXR �jW��X����Z�=,--]�,v9�Ϫ������FZi��S�kԕ������i��8x�*�FOhb;o-�荎���f��	��n�7�X�Fu��,])J�)V��i:��{ї1��|�}:��f��$ <a:�͌n��h�Ff�"����~�L����d�+���`���@���T7��|H=7��ֹ��@����`���v��~&��{���Ily�7hSGً�b?K�u*7�js��b��ʷ��LMm�?�WP�'�����`���\�H�Rǟ�|x���69�J�a�E���u:��1��Rq�g}f��xy�F��ӷ������<W�����JJJ P8o#[�D���W:�=]j[H4���˫��
$��������:ӏ����s#�1P��!���/�6��y�X��D��u=��_���IUu�Zf��?�����F��z��X$2ڼ��쨸%b@^��V����*ւ3x���nP��Ou:�
���[�RǨjh��yN��@��Z���߳,��X���c;���*�?�:Ψ������*�������3F$sq���F&�@t�kfM(�*�s_�m0�ݏ�`���s��jȔ^���R�JEm?[����8���7��j�"��6,��!"�6ߊ�.�Gg���_�ڂ������kX� ii�$w�b������"OfpWW���&�}S��Q����,�������H����R9�r!�t�,Q�bH�!:�����K�M��4Īz�e����7������\G;��ҪY�B/�#p����jq!*-�z����΋H8�z3D��Xu���Q�+.޿n��X��
�°v��2hG���2��:6GT�$��n�����	�?;��r?F�1s�>� �Pr��9���V��'n*� �*����B��į�Ƴ~v��I��N��d��}�� ����G�m�L�x�* O����yI��⃃�$q?�1�}dP��F7,�=2��M5��BHKKwTG�,'�X*_*�qŸ��1��ҟ3/�S^޹�BJ���փb�'Rֲ[q�ס�Ii"���IjY�������@��2)g����mR��i���V�3�)F���ƿŢ?����,�8]�V��}����_D��[��n(����
W�\Q56������]�Z���� �*�F��&Ʉ�Hj�A�՚͞�p��>�ȵ�-|�U���>�R����NV�x��MC��ڳ0-~B\��Q3�5�a�3����-���O4��������^�"��g�* 8��{o��:P9������9�'��P0�>��n���7��8�I�[���5���W%vd� ��Y*�]�d�p�ٗ�R$�;=lr�1�c�3��d�&�	St!�@�/J[�#8���N�#��aSX���R�1�4"%$����OM^~��%���(Ak��H�R�=s�,�B��'���U��
RT�}y@�)h+�3�%�G���ְ�Cw�R��H���uy��؟���+�%��F^�y�;���:82ZVB�����{�}�M�q�}����{X��ֽ%�����ǋ�~��C^Z�݃��j<��	L��$��D:eV�}ܶ�5�E J"�I�A�w�GG�	����|��̌ ��:���)R�ݳ*jB`��G��!�<�Yt[2���S�i���`'/x���Ȳ�����Y�6#�FD\H�O�DO��r	=��Ron�J(:���l/^�fXXs?��%�mK��>-�P=aa
��)
/�g\��=��猈��X����)�̥�T_3��{{;�j�C+�-�QD�����*bɘ{W��� ʦ��V,�:�{1ϛ:��`s<!T0�N��{���A���¢W�����2̤g�E�$&���� �;���F���nX�F�'�7�8���y+�{`o��?0��Ŧ7�����uMG|�/2�NǾ/!y������F��Gg�, `4��(e�Ȯ���~g��͛;�U����6��<Ɵl:���T֑���S��H�x�9n�iX��JB�ɵ�E#R����}[! �v�--�ka�,�AJ\@��4$�C�����F����`QN��M���{���}11I��XQ5�Ð�^i W@�����:�����	��?�ݺn�a���rcnsӢ;:v��4����� #u:|�Y�H��I:Ea�7�5�K�|9��?(�2���,1J�J�#sy��,�@;i���g����6a7��<)N��bc��m��|A1׽�=��%0��,����qS�
;f4��:(����Q��=7b�M��M�s��ْ�J�r�g�6�y�=��R�6W}�ً_�זҎ��j�g�rr��{��AY�n#�N��wfj+�xn�1w]G�*�])�%O2饙�Z'�#��RO�_K,�?Ο����Z0yJ�3`�`6a����R���8&S� �T	�1��מ$�؉+	g!"���Az;�{[:��
׊ .�.�djsK�b�O��I<�6w�e�1&-q1�|.������"��E>G�g'�5�^��]�����q.M�mA� 
ԕ�'�O����s���>�2|����0pq���^&��(�����9��T�Qq_�V���ͳZ^�W���(�]����lu_{���T9���mC:��� LP�F>��ԸH��W����RP�i�RJ�^�tD�����o`7��0�Ŷ�`���i+�\٦�Ŗ����DT�"J�#��g�v
��~
FЬ��SO�7���i:z�'�����σn �-Q�L�/�UX�b�M>I�)F�m׎L�@)���N��{��(m�=�7��0������ �����{[���^�!����8����1�u���Z�!�J��׵�w�&�.bfo�:��ڂ����jĕH�x�td_�
�����\C}i`�D�Z
˘#n,��w�|+PE�"W��N�R�>a�o�:c ys�J��	����M��/A/ ���6�p�0JZ�>��H?	a,���hGy��N�c9B����W����>��QSˎ�ᘖ'�k�r�"��b ��Ɍf�E�޷`g�O�*�>z�LN؛RIhOY�f8޼=_%��V�����gw�<l1IÇA���#�=4l T�K�3)x̲�N��x���[�;�� 4w�v��Pg�$���:S��8�֍�ⲴB,�)�_K�Ư ]W��>/߭���aT�l��h{�9��]�|s�5��Զ�������Q�D��a2�}2�{#�8��a���Jwf��t�Xa̵c��X]Yi0x����M􈾰"���L�~��!X=��H���>ث��8���NO׎�iG��ζ�s��lz�~t��hO�q�x�dro�/#��c�|��v,vҋ�t�"�)��~�ˡ�co�~;@3M�"�2�pp]��wg�Z~]�[fs�m@�%S��Α�^� ;�p��ώ�7������H4]����O�*��OL���GKs�zp�PΦ��r_�����ѿ�H���h9����t;�ݏ�5�֚5��?N��Z,,�;�Y����`�A��`Tb��s���P(rr�H^ӹ��'��G���Ҍ����������!��	����|��}��[�Ǽ�ϭ���yr��/��S�g�hٙ���G��,D����x97D�r���9�h�R@����ʶ���D���d*�A���P�	�Ԫ�Ō;�J��NX��Jk��.h��Ѹ��G�4^�[SEWhK�ۨ�E�����Z��C���	jg��% ��46[�����="�(%M";�,��t�{��6�%��ԛ�
�Z�����SIS�� ;1u~n��L������|���v|�qYHmjL����c�yۥ�85�X���Ό�ω_��ƕ]�K����E��b�9B@��It�`�!J�3+�Z�٪���:��vr{=2�[_�}�gjUE&v��7=���`ԯ��Sw���m����5:��2�syQ`�@	.��چ�	�5b�S���|,.���dRn8�t����7T2�"�}lKM"�j�wR8h�ݜ�v��w�f|7������
�v�M� q�!C�ȦT�;G$�͞,�V6�g�xVV�B�����i��k�͡����- �p��=B�Q��mG�>�S�F���8-t=������q������Fjq�B&����=|�X{B��B;��C�(�v��L���]����Px�������R�/�:Bh��N���4��	B���|0`�<���-��p0����C��T���gU�_Y�8�T�[�GM��	� �q�5��R��e3�f�p�r0��K4�Mҝi��B�p(N#�6+���?:3J.���'�m�&x�`p"�`VW%�,n&oຑ&h��2��_v� ���sOXv~a�G�����P:26��[�c��>_��aQ�]��_2��T�`�iS �O�x�����ҥ�Xuf��[�뙢u�k�@@þ�����χ=��)S�Į��N��>z�ZQP$-7}���Hu�hB)v���_]C� �Hi.7��/T.�����7
*��{cWυ;w0�'����<��+�R�Z����+�=�7����Q"|'� )�Y��O�(�2М��3}����-ο{��N]'�=C���)�.H$m}��5U��k�N��G붎�W#:>Ɍ��~_��͸xo/�ģd� k�bu�F��&T��Os�2Q ��r���`тO���������
�6_�2K�bK�=nu�2���S�)�̣�P�N;���q��Tf��f��Ju57=�=�Z*  ���% �:8Hae<;�gt�&�������Ӯ�m��-2�����K�꣭"�Ƅ\�~�=)��N����+
��kt��� g�������_��֥�рI��H����V��t�c[���XQ��{>�r��so���"N{���A�~��`sZ�Gc���9+'��Wq{�p˵��⪤�l٫�?u����Rlp���R-�WC��.���gD�BnĲA!.��8"�ԶP��紜�c�
��k:L=�m2p
v#!�~�Gb�@0pਣ��9m)X����Խ��}Z�'7~eC�XD��N`�f�J�R�bRե�����d[�=�cj�<��sJ-Z p0m���[U��:��>5��Fn(~���s����(b�/�7�Yv�����ʆN�7}dŀ ��'��&��t1���́{��7�O`���ut��ć�ڤ�⯕���$��$��e�[�6Q�C 7v��h#�YR����C�X���J�^��[)'~��`q�閦�����$��qI�� �x��O6�l��ޞ��&����������$$P׭�rT�A���������£tܘ�OTٰ�h]�SQX�h_�k+�ŅJw%g��S��LAFe��j�L��r���;2+��_��������S[?�e�Jkz���z'� hd������?Ƅ	��6Oe�i�uVy����p�KPVZ:������5IB�(5�ٹ��X�]�Q,��O��82YC-�k�R�&�dɲ>�N2X�{��/eq�I��&��b�ٙ�ڮ����d��p/��)��1��Ȏ5���]j���������'pW�#�~�)m'��]s��QLg2$��E[D�Ţc�. ��'4�<CП~�d��� �$0e����%�P���.���������Z�4U�� v�l�P��y��
�H��zr����F���\��HM��������7����F@L^G𗋙���B�q��f���x]��1ѷ�������|*"%�	]�6�	�K�"�G�:n�$.m0F$�ߕ�4�r��'��a�����<ap	��M���B�>����!���n����g��om���6�o��c�=�u��ZХ���vR��m}��:���J�6��z{gG��
/r��IК�C��;�܇G'_��H]z:֑��}�"it�fi���w�)�=c7(K��>���E%�jLU�)j''��Lw:ĭ��`06f��A/����N����V�)���)+�-�$7LoK��>�~a�BWs�=zR����✱i�
Qy����[�u�u�j�U�+��ؘ����j�|?�T�p�}_"��~}���yqY�O5;썍G�_ŷ�Z�y��˥C�"���Љ\���&L�jXeǼ��� Z�e��O%��ً�)���4]M܄ogz��2��*��B^F�Q�GU���f&>y.;�F*nM=��8*j���\b��ܸ�`}�[%��M�K��*�����1m�0m��O��ѓ���;�:A����g9�����d:��G�� r�`�����]�[�4��U�������ħ.=>%*�R|lF�c2k�I1e(�`�Øۡ,O����W7��Kc+��BK�@6|�����c���d���o�Ag����^ǹ�y_=Q�Α�m�)��eC�=��rx��V@��'Y�����=GW���,]�/�Ƙ)�����t]�`;��<_��|��_G�h��B[=�/��8�y�h��ܢ��W�uq��<�R�*�}���c�$+�g�͸V�0�@�N�shDau\�6�8�
�?#fD���0ߋ�6�Rs��H�D΅*�T��G¼4��s���rBZ���ߍ)N�Q�ׇ�ifq�35Z(g(S�K�LT:p�P<��wh���ܨ������҅��,��{�s�������:�|b��YxOJG�l^���Pl'#�}�(�t�J_!n6�-��Қ]�0���Ⱥ`y�x��v�^����ʗm+�.�1b�2����������Q��K��ڋ?�j![?R���ew�/���s�q�,�e��-hZs�s~�*�t-��1�Â���O=�T{�|���7ښ���sA�7U�G�7y9�����:��}�}��8�f��3<j��ZE5���~-N��w�����&��$#s,[�,W�d��9!�/�7݊��&E�a��JM�Mff��V�q��R�X���骩Ň� ��\1O�Ǆ[nI�g��y�L�[��X�Y!��+����Ww�����tT��������u��s�Q��x��u�T��A4H�3�Y�(��=��o%l����_����<%�.nC����w��h"�B����t��۫�dl��\e�f��d�����ܙ�����sZ�=0����[�����|o2>T0�M��;��&�����M��F�<���[�,�7�K��Vo�U�2�|�]����l-֛��BP{�����ׅ��9y����uܺ���6wfz�)n�efw�Ruzmơ�i�Vj�t�` R�jd�~�:a��D>���O	�ͮ�3���Z�c�o�������ش�%ZD�!�y65�(ҙf;�,��r�����J��Ρ"k_^�k���F���u��빋~��s}�M�"q��r��	���M��-ɏTފ��Kb�\��IU!�������O�G�z_�����J�Z�V�!S��	`r8�r�t���&��>���Q�ⵆ1;H7�@��*�w��S?Ǩ�����I"{:����Uu�f1}�R�tM�j=�S3�Fh����yi�RC���K�};Aoܺ<|!����
��N���p)#%�ӰS|�IpפU'�z�;]�I���f�XEo���f���W��!N����$���m�;2q�,�!|o\z_0��k�>��c�tLR�����̠�U���E�xawi`~S����T�Db��X�]�Ӽ	Y��v��L�:wX���mw-���dɱCNQ�� 4�(��h�.�ޠL�W���O���z�+R�u����ǖN.!��"-����"l2�e�5����B��E����ۼ�k��-�G��+ۡ��9�:2+�3Sc��j�*�)�ft?ģq�|Ol�[2�on��߂���x�@�K4<��1��=z�l2~''��
����@�J����cv�o*^��7~��ϻ�8K=RE��z�+(�XN\�@�ȷD�^�]��E�O$�8χ��I���;@D���y�����4������u�e�8�8�xꕯ�u5��\����Z�1��q���\�-��Y`�-eZ2(U}����]$��~lU��ܑ���7�wN�F;�9�p�7L]���<=�l��3�J�8Y��Y%�)_@�v�'Ox�?x�b��{����c����P�t$��]���ꜚ��T\?kI��]�zv�m�E�<��T�P8�dd&�^r�` �χ���2M���6Ui���[�n���R6�e�ܓ�e�Þ�A��'�L	M���$h��m��l�D�_��;Z�q���\ȳ�͍g���A3ߏ|6��A��Oğ3_�;�n��IcT��a�k�:�C�a?���YxkY�����.����Է��*/����P,��p�w�n���TBq*�~�ˤ7��c���C�Zf)�)r�����g����i���{!��a{�Ÿl���E�v͕)��~8����Q6��7��>��j��IO�}�(��u��|�Q��wo�Qu �(��xu��lvi���2���������q/BϕV�O�#�� R-S3C+H�~�U	�X���3QT#��Z�P���������>�"؞h��V����n �R���$�[�����:�����92���yC"M��%�9C9U�rC ��ڹ��a�9�4�lyk� N�qB6W�	�'�E�x޹zMn���P�B�*+�k�ە�P$�(�i���2�>5iN��ԟ�"�t�9U���u�"��r v\�G�(���[cv��w,R\!N'�z]{� #ڸ�n}�V�Q�33��f�����S�.elќo2>`�e�����ə����RTh��Y#3���
 g@���D�l
�55���s�"j��(�t�՟��4�ҵ�����V���e��MIyZ|�SSn��>	H8��2�� �z��sv5^`+����E�}S.]��N8{��Tǖۃ17m&�1��Ѐ��������}����+i�d!t���A�[���?v����[���,�x>�w�x�OOƪ��|t���b@yRrI6�~�c��n�M��- W=��� �ql\y>�T(�X���R��zZUV|zAY֮D{�E-g�*� g%
2_9|�"MB1`�'87ѓ��:���:bn5�Ftճ.%���f���Dd(�m1��^a^S�F���?�a6���i���z���X7-_wo?�2Ά���<@���]����y������W�b@���s��K�+�@U`[�c�D��,P��z��&%L-o�>6Z�8}����Yf�����7|�|`K���Y ��o�1���Qr�9�/b�2<�۲?��_��rQTn��d�o��3��`���ӌ�ƲJdQ �n�(y�؄�?9���V�y8��RiCz>�#�3�����?����%Z�#���8��3*��i
xm�zz�P��� �z�I�j���Wj	-1$*+V~�����4���td�鸺�t����1�V��eX�@��^e�t��@1LX̨[~{�O�q���p�0Bw]�����IoojT�B�ғ��B~�?\�\����q�뫔�C�j���'Q�M���1�;x}��w瓹��e/dEռ�T��i��D�W+w�P����µ��־B���,m�^�McEf>ÏG/����� �LjX�@ؓ���	ݚ~���5����74R"��K�ȕ;ǚ�ɞ�һ:�7܀��ܲ����}�h�S������s��ϱ(;��\R��̉Afi7�(������W��(�D�5<����Ss�0����ׅL��е���q�a�����7&�.T�]z�h �p�o�-�j������D,�7��(W�JΟ�c��q�]��*�z${z���؆���DI!Sۀ�䂣��i~f��7
�K�=�}r�����e�9�P�'%�R�Yke�ZvCg&�4.�-�\����������9x�J�e�Y����q@aV� �+!T[�TX�e+ߜ̯}���2K* �����ȟ�UtO�8��ת��T��Z�{Cwé�F�.�zj�b� �y�����G����v��������H��u�-���/B4��|�4|�G���B�+0C����vQ6����ܗe`Wy���2t��?�"���ѫ��,0�|gz*�^��p�D�`r�nJ88���:�` �T�~lu��L�[B�1�D�!ܪ�聽��������3v�R��+~��4��9�;?�3+]&x����
2j@> 
:�~S 9���rC��n�K�q�	#9�S9n��t�XT0Sm7�%��I�i�<�y|��$��H�)��b���Xh�0�ve���cO�a��g��#&5!�6M����k4��Mo[�$E8{7���AӢҏ��3_h��H���s|@��[u��@�����Pj�K�P��Gi�60�}k,�k`�pϮ~{_�����{�7�U!&6��գ�' ^���%'�&������#9`au���Y���$Ǜq����o��4�?'(�L6^�Q�sa���A����3�d��������[�Y�To�,�`׆&���ũ0�2S~����B�=E �{���>�"|����IOh��,om����|x��l.��uG��t�R9S���N��
i
�%�
K<�D�ߡ����RQJϷ�i���3�=Fv���'��?v�̣�Ŭ��y�\��u{�>�(u���l|�+��P`|hݨ9:���mg��E<l��� ��kM�%',%�ׇ�By^r��-L�%���j�dʅ9�?�7���'����qrC=�+)���J���+���N۰@sE�F�/�<�ƗF�[}�����Y��W78e���`��T��-�,��6�&�󺺻 	eKT����U�ކ��N7.t>N�l+*Y��q�1V��$d靰�;���i/k0�����[l^D���C���۠A�gN�_�F�e��Z�h�a��p�T!�e�	��E�D�UF?��&�B5�XPє2
����8�k��?:�@w%{L��W75�@��q��?��w�\ 4��Jǂ�-yU���#����	���\1��"q���d����2-� [Q_cL�2u{[�t�����Dq�$�q$A2�!��vOO�r�gn�L���������5��������cŃR=�F����?��I�ī4�B�c ^��4�A� Ei���>��)�Қ퐖QQ���W0ƷZ�������M������� f�h[b��m%����w�M�k������}zk�8��[I��k���W�c�r�2l@�F�q��w/8v�������X&�`�@���3q'��9ҍ������bV��l��O��oё܈},qP�f�!�H0��\��ߦ-w�Fh�)��Ҩ\��F0�D �g3.3�.F�O{pyp}�	СʈK�#�~Ы˒s���vr9ic���Q�>פ�f+���9�Ԫ����b��br ���<;<C=�a\#�u��|${�5ɽ��B�AM�.��J���+ufz�\�t�u0�~�"�>��<_m�^j�g�2�ؑ�V �V�4�䗒�k���Ȏ�sPjzZ���%P�ގh�
��j�v����{|/�w۩����I���k�ۄ�����e5  .�s?���7�7����L�`�E�E)�I��r��?2򓥥^���.�\�ξp��x��FO����o0~��ܛ��[1��t�#1�Bؑj5 z����V����2.��e��=���i��.��%ߟ�7.@��RN����(E8�.�+&"r�r�zDg��u�Nl$��,�"L�Ƶ�� �i�k/��1�=2฼�T��O��ڃ��%|z�J9���a�K��7�Ζ�f��gh���7�Mí(��|��A.o���8%��u�EMN^#d�ϣ���=:��6ۅ��6;��p�P�n?���G��S��π��6U�9�P�8h�� ����3&ʧ_��lS��c�*�܍��;�]���	���No<8���3�1��l<�_�z����C������A�69�8[�@����HΪEŪ��ӡ��	�_�Ϭ�>u�sg��[�*@w�v?��*�^������E}"�6md\ɓ��=t�^�B:��=S�gvl�#c}-�^1���@�����W�J���jt�Zq��U��f_��s�画#.�l�V��G*���?UC��z0d��ǖb�
���&����w�H���u����pכ�~�o���	�q]�,�麲��f2�T|����.����غs����-���*����������m���U���*i�Ο���LD��T������ƌᬐ>�>�q7Ap�(�A�P�/����5p|9��o]8��eo7����SK`OI�1S(5��v����1��2���1D�4����� �.�}|:�_c�e�_�H7����DS�� ����2�������'����pՅ=�ٷW(y߼,5}�ܴ#l��cӄ������<+��~k�>�w����[���&�F����'3�����	y��`��&�f`�P	0D��?4�]
۸��eV=��uWOψ��4cu��X���~�NeނB��h`����� A��ϩ��j*i���x);�;�G�=��OD=P���uk�{�����Ï�;B� $��n���ҍ�ޖ)���G����o�@-[�A�r�����A�X{=%}����1����ܧ�%~~����3ݞ�B�V@� ��Y9��Z���[��y�#Ȩ����N��Z�4�s�"�n�T,�J���6����| %�3?���3��6$'����[�?29���B;1�&�j�C\�Ř�eu���w	;�6uJW(�}t�Do�`��آ�@}mN�BSq#���h�W��������N���/�\Ɋ���&}�,
J�F�5�-���9e�ۃ�/%%�ڴ����u������r�dM��/��m�ɭ�o�c���N�Ų9���+s+� ��{�Z��e��	)������p�v6��񁘦i{�?�XaIy�||||�!Atӯ *�vR�{Un��Fb�j���%������ /*�@+��Q��An�V&��؟���MT��&��"dk���XE�����{�a��/�����.�Z��TؠS��,ڔUb����ӜN��2�ku�:ES�̗׭5.+jOӕ%+�9,����3O4fOv������n]X�������U�w{���nt2ڬ�9	�0"@X�b��Ւ
~��W����6�!���3��O�ه��v�{�k�8����8�5����:�^99\G~�r㦮����S�2$�W7d�� ?�{�ӈ��?�O�H���5��,��!�*��ھ>*b!�((�t+
�4H��t���) !���]C����C�4CJ�P߽�}�7k�d-�{��g�o�i�,)-��ӄm�6V�Gr��ű�1�\ץ����ˆ��t�	9\.-� |2�����/J��?Q�d�#�����F��%��PJI,]<<&�x��[��-�r�������<��T!)�/M,u���	&Su	�6�QQII	f���6{�Nɉ�ބS!!������WU������9sٙ	K�kT�b�#˻��?{��o���Ԝ�ڌ���2?�
�	U�W������å��=��:�����sLn L�['����c��ʋ�x��"t�W�$CG�1����K�t��d��ڋ�ل��\�c�t�YL򠨐\�G�e�V��� Ҥ7�����T�ׯ_�l�h��#�ֺř��#���w��]c�� ��wV�����b^�xKP�j��pX$�����a	X�-�&{�uttȫ������
�{�U�.��Ω�B.�:W?��� )�U�;�LH�����n������"�D.o,�Ǻ�K��b��x����m�������}�a4r���e�8���Q�3_����#Li�c���=�GA��ʤ�Ä���D������g��8y� T�mVy��A7k�,�h�H�@�\��8��-�O���:%�iJ�KY���?Rz�\R�|�������o���A�F^OO#�?l��l�?'���SW�"�B�����{kj��8?�Қ���>	$K8�0�ak�AW�?T�(���@��
שj��53�<����"�����ic*:�˘h7����5ȌX��tu#��q�g� ��[c�v�kGB�э�+ Ϯ�� `7�m (7dTPR�\ޡeb��t�c���V��m��~�
�j�[�������������/�C|-��F�{0�
hl�B���I7͝�o�J�G���Փ�<�t�:�d���d�C��F���E�W�с3`� ���e"��R��


FM�w����\��&4�{� ������(��	G�9��7Y�L�9X��+�;ou�)Z�g��	��c����b|<P2��f����r��랍]�ȃc�q\2l�����4~PE	�!���[�>���:U�g��ʩU�8��־���yю�N]9�)��%%�bS��B��L�bؖ�O�f6�#�5��]A����  ��_
m%8�?V�Ee�R�K�&s@�_����Zk�b��Y��e���|�� ���%Ă�Ab�Y�k��(��"���z��66#X�.�I�j�D����A�V�t;/]e��jf 2��W�O�X1���g4����BC�?9X�L���_��7�A���;j��}�V��hpQ�,��4���aؘ�����JL�7񦚈W/�|�19��p��W�G��E�se�sE�z/bSJ�I�UrdH5ૻ"�����������!UJK���Y�>��$%�dʒ��!Zsω��Yc!}q�F�&�4�2�i��PI}�G�l�� �)����.W�Gݙa�)�$���U�E<�gv�|�k����x�����k6㷽^�c�,1ZIz@��u�����?���I�(��M�ҍ�q0&XA�|'�9lrA�{A�S�ESf��u�rʞ٦k�����9/(h:$K;���4�v|�Ǧ�� j�n��j�~pϮ�v�Nx(��P�NjǴ����7���dH���ތc���eXD���a���%`>ǈ&g�\�LI�V�\E�N($�}K%�_�ve����/��Y�}�1p�w3䤸(�N��qW��^��j��o�p̌���R�8_�[� ���!\��Y�x6F9��Ny���Ck��ё2mq��m�����0���눿��n�װ�����7&{e[#��}m\!�}|�l|��0��8�ɘ��)߾}�<�oZ�9����Om� `a-�H'���h	��ڰ�w�b[�宅�)T��P<����-6��x���o����pJ�C�S�5u�=Z�1��Y�cS�b)~A��I�lR2Q�t��(L�s�1�n]}x> ��{R#���Nq���_	�N���Iå���-�R� ���@��4�ZmQ���o��]�^���L������gP�	�I�������g�N��4��f�ډ�F�YhK��‿��|aE�5	�W��[�L>-g��1p1v����@���,@:��$�ϡ���i<��N*@����Xn{����WyUb^�%��'�k����T�����w���q�1e.(SӃ��>�V#��m�FX� ����( ��ץ�����k�3���0�l�+y��N��Ǽ!RB���2$yt��&W�cQ�KRv@��P�t婤����d����!��f�q+Y�/�f�j�?�[a�r�|ߢ����e_7��;�Ⱥ�����l���zx��>��c��<�����,���Q��X��x���[�P�f�L�f*�ƈ�Hjo�p�Ou�??�m).�@�ڻ�ʥ9�i�Ke�쉧�,���OKG�oVU	�6��2����@[�9� ��M4�WR1
ݺ��㟔E���䑪�7�&��.��ifw��^sK&؃:�v���F�f��5G��8t�7���$�(d�w�\EBİ��8N��`}�U��&����]�o	�~6�9R�a)�B�1���6@�;���K�\�;h�'D!�ҏS�\�y�Vm\��r� >���N��BY߫��V<��e6,ُ�t���bc�O�]pDiY��Sѥ�`uBL��9s'��z���|�W�Z��dE S-\����`.z7'q���$T�n�������kre�S�C�,���a"��|NmIrc� 7�v���QF�J���+�4�L��~)]ŗ��$;��9�qX��ɤ٢#�r�� 8���$�\Y@�x�� � x�����6�����j�IJ������S)��o��4&؂��;�����-D���,�OF�[x�dd���)4��α��$X� �@<�Dv��,3��V{��nػ�`��V��ɉj�\��s�\ik�r��n�L<��<���NI0���%_���~i�KC�3۸1�ы�����l��Lށ��Y�U��Ԙh����ޤ�tr��&�:'Sg��1�-��Ҝ0�MKή�7��t����d��X_1=����9��[h�a|�MYW	�S"�2Dn/�Ǜ9�2�+��2��ItD�����%�a�9�u����p�I�y3J�0�<��*�.N�|�9i��}��Y{Ԅ�@�yZ��:X�Y��n��e�-�z3*
�fxg�����:��0��	���yq�l����(ꍏ'� �p�$��2�g-�Ӄ[�km��0��$+6��)?�;u��b�"��?+�D��D��K~6y�B�Y��ȑ�W���cW�pm�`��>c�A��7EQ����-���f�����$��6Q�`
�� �H;y23(by�RLǈ}M�}����4%b��O�N͙E9��e#�%N>�e25`!a�Y��[��x���:�b
���5܍��|��=�"�[!^��{$�����	���zҨ�W���#����wR��(�X6mֲU�����{����~�P�1�r��{�����I$P�(�8���n@����2���9���T��O� s�m7���Erp������Bӈ�ΰ�&e��!�C �m�R�%��7'�Ʋ!T,k���v� �3�¤����ӏ<jLآ�[.�o�A~M��	�0R��8x�&� �f�P�k,��Ǖ~�X+��(�x�w��j�2�,{ӊ/����	�]�O�<��fШV�i Ɨj^0Z�5��a!�w�"��G]j�������O���BT�z;
�R�;8dU%����ZX�KBG�b��
�ȭ&�s���|��;D�櫤�/:�R.`��oQ��"
 h��>/3���~[_qg��Lz���E6pYI��(��$���kvF]R���=�!
�Y�uhΧ�����ۧF�8�C=u�S��Aۙ��)�~ݒ�3jW�γ�"箸�.����թM��l'���dn$�A�6�7��x�,��ߔx�c�Wn�esJǆ�q�Q�U84k�)0�����5�z��xy٢� u�&yו
�O:/�U2����)4\�Q:A�qJ�����
%c�$lt��<�v��
Q�{�����sBJ�._���N1�ϙL}��|�S�{Kv�K�O��;o��L�S��ce�W�v=�*�WZ�x���0�e�����u/���]ƍgf3Tl��q��JГ"������ |+�J�����G=�D�J��]Ж����rQ�N���Ǫ�1��\"?�2�۷s5����`�(���C�<\�s����Gtk�G6W	��S�މ��/1^�zn�T�9{�OJ�; ��播�����[%;�J~%�H�������_�8�?���O/[���/Č���};����yd;Dݺ|m�V��s_}Q/ J�$o���FL����v�u��Hߦ�6=��͞xr�q�i�%��^w���qg-� *�J��#m�R��
]�RZm5/u��ƍa�"��\�69��so �v��-�z#���FCArb���ˡ�A2�u�v�Y�lʫ)��q��.��t\jH(��9��B��̒��Fp!�ʗ��>���y�)i�IՉ�=�J�(jW�<k��y�x~�C�A o�#FUS�i���H�w&[m%^Otp: )1���=6(yS��>�SO�*4�f;v�Xa<�
�j%wu  (|����!�/�mY��av�b��-4���a�E?��	�3�V 3�+|s=���o��S����8�y>��u��?��'2�+��;?c0����>�*�ǝo��M���$4-1�_�e�·���W��c"ް�*4�5�Ù��x*>�F�x���C�?�9�c�k �|�2��s�t���-^_3U���"������`K��'Y1Sr�󛞌�7ӒΩ���a��-$���T<�'C�Y,7uH{Ow(Z}%���L��u���d��s%�%���k�7/��ci4M���C�&?��k�D�V�}"�'�^Ae,b|�n��o���;p_>8:�\$��d�H�Bߐ��Ҝ/�=unD���V9�x��qu<.���l0��/!��TQN���*�Tn�#�ψ#d-aɜ(�N�K���N	�~|�����*R<"�N�OW�q�~s1/�\���(f�qX�&��X�=���O��ݝ��K�"'.�K���G��7wt�Cm��u�ׄvl��YXXX��7����nQ`y�$�05���� �ɑ��:��U�䱙Gl^������5�d�X�7�V�&�3 �uW�b/�^�6J�G��.Jp��G�cL��@<ϴ��o�ב{��S���ף}���U�M�����zg.u%��=�f ĩV�Q";T�12."T�o.k|���Kc-�"ԭ=0���*"�!G��+�ǯxx�K�^{�e�k{$�8~=������������ܕ��)K�&�z��+o�\(�}���,��S3灁�A�޼���8��jc����j�3λ���3� G���9�]21Ͳ�KpX���E� �q�:��Lҿ!:a�>.ǠDB��1.�aP yv����ʀ�y�~l�]f���������O������`uJ��f��^���˻	�/O"��}��ƻ�Qi��V�ջ�.�68{�%�8��-*�"+�\�,+:`�vS���8�dN�(ބIv�)LI��9���'^���~����@�� �Аgs��t{N��x�{�U�]��5_@�����f�$��E������R�z�-��Q���֥�ƺ�f�;�Ā�In�B=W�#͛��rpm�����ȇ'�dp�Ro��5�v��z�P�5G<��^|a6�W��׺�~���E>�Y4��1U� p��VeU�bY6���
��to��iU��
��s�����@_�9�I�9!LE�$)ve>��&v����˨���p*	�$�� ��x-�n+�@��݊���Y�Vx����/���}��Q�'nO�l�7��jG.�h�)?5��V"��ƣ�|2�x�����_p�N�ȓ���ol���~�3Q�#�2yp���:CN�% EN����7E&��+��f�fP�r�Y�+���_��"C.��T�T�+̡�/?�2�Bk���S�פ��pr�h�:6y�ytt����H�����eء����D�ź*�3��_%�+!����4�aA�o�&�
c}<x~q�qP��p���}�/�~YfbTi�m���~���qR���,ߵ.n�����[��ѱD�]4��)�ٞ<N()Y�[i�yc�P,#�k���C��cr�nI��� Z�*�N�C���;ȡ+�緈ZZ�UY֜���
��!\�R�����P���.cS�~?*0Vn2��_9�LDp3��'��H�QGw����7�H�6���)|���7L��ll45�mqQ)��gdy(��H��N�Fp���&�R��!�7$n��H@��X�L�S֔���!7�Oo������!�?�o�o�c3�������d��3����a��`?}���e��>�=66x���H�p�?{�HK�����l��������Љ�ZX8�{̢�U�������S33���gQp��d�G��z�ផ�ryv�#�z|�OP�^'�s��o��;m{ݘS��.c8���ɢ'��mć0��hNB,��U2��*^!W�d����):U��ED�,!h��}��.ԡFZ��T#�ñݏRV��L��u�Y�yëJr8cZ�V�e�45���B���*��S�9wc�L����"a4թ�t����p:������5;#�߽".�|qw�UZ#�&iYvS�.����l)m{��Y������_�b�^Φ.�L��r꾃�ѿtΊ���]�R%ا�CGO�)�姨+�)+g�uFа��`��m��Lq8�w#��I$b��Չ;%���+�{ꃛF�w�a���J�����/����X��Ka�������R�11��'t#���(g��� ����?+�b�D��������/��#Ww�ɞ��1}ݯ����@q�֚0��L��oI���N���EF�U���b��l�b{��zm�!d�w�Y9��Q�*��09���턜�z���?��e���Ӱ�{�x��w�f�7��l�ě\5�n\*e��\�VC=t�ed|drA?-S |ٰT42�@��7������|�ω���2Fv�d�uL�捂�g��dvaAd��G�.}�l`��+	���vi5=�5½|���B�է,m��td����^�%�/S�ꨕ�w�%�u�@Q9�D��@^�Y�N�)��x&{��Ң�U6�1��}�3Ipd$^�5�Ϊeo�1��h5���INJJJh9Zi!��s����;��]�p�4"v��<@���[����z+�8auf�.���j�9�;ZK��Iy�^5�c��t7�zh3��;� 2U�+���}꣐��=�;�б�,���)7F���j|�H�Q�q��\�̾b�y0dҺ��h����}|�$�`,������b/���(���(��4�Yr>���'טkvK��+gn���ǝSN]�h����^Y����.�q˗G��\�$%%�^���p$��TY��5���_�GY6��X�<=���{���O"�� �51����lш���r��7jrI� d4�x2�FX�Iq�[��$}�)L��x~+��,�o��Q�O�t(���������`��Y�϶�t����m|�9'&�4��Th�3�g6�
�z�br��*g,!6������^y�=��c�/XU�kh�sc�cYZ^��{��#z%G��.���ԓ�Dn��zG'ώ�*�8�]�4��B�=��jF�o�6���EqL��,���\�OINV%,|Nd�b�;���D��R��i�A�֭Ӵ�x�)~m��k
8������J�~��������G�2þg�v�.�s�J�jp?��־dЬ�3��ͷ/PX�2��wٹ�t&��o�4�A�#$k�F�)(�W�Ŧ�t��Wl�;Hֿu\�����v,�Ȅ�Z�ڐ���Ͻ��������w��(]��#	a�΢9��nL�g�,O�R
�U~��^|k�^Y����wcvn��Z����Z���R�V��q�ꧬ|�?Ku���zz��1�}��`?e�|��:NK���N�gAX�cwm�_�jNmQ�"9�i��z<���,3>�鯬98��"9��;8�x���ĕ3H�۟^���XASM�*6z�;ȍD<���&ώ.��v�K�F|6���nF1�C�A�}�A�+���7�p����T��UIX�6��.Q��.��a�g����r8��.+��nR�1�t��F|J*ۻ�sq��1<c�L"lW���PW��677ˬ�:�"F)� +�&��P��4E��k�+��u�J�$#T���U�K24�e cQ�v���U�]��7����!��Rj���� R����P�9P:GM����Ɨ�}	]�,V�2<����V[�g'7�6�7�j��ؗ�g�1�+:�H�v��+&!�L�~����=�ͤ�Q�r��g̗��j��������E9n��Z�P����8!���=��t4�_^u���"��TK�iU)ZsPB��d�@	�$�\F�KX��f[�"?�S�阱����T��:�3��z��|أ��	�h�������m�+���y@Ġ�Ln�%�����YP[[�U�&'�
��}Bdu���n�V�tj�XʥU��h��6d���,���8�u��Yz��Nu%�9,��cϢ�v�P�<�]�;3�6K��?�N�O���G=_!�6"o
S?�:B�Y��K��qq�0BR���c�� '��ӳ"�$��R� ��N��HKZ5L�K)!v,��J:�K�V5����*d�.�ua�8��|���CC-���B��������
��-� &wY��*\ǳE��~o"��ǰvw���O����w�k�g�-Kv��&9p�]���&����:�f�]Ч\��v\0����⋩�I�1��Մboԝ����ۋ�A�f�>Mɟ��1��GDFf$8P.��6V=Rj �?�fv{�*��7E�S��7<�>���%���I�_;�����-��@&Ջ����՚��V���a��O����6qo���Xq�ԫ�RW�|8Z��e~�NBpP�T���	#?�������e*��������TJ�Nv
S+ ��a�4�*�=��촯�l�Y� [�4��j|�/x�r��_:���ȸ}ÿ$�lѧ%�^� &���pS�G�t!Ŕ��C����@�B���A}1"��-+�g���Jpx���jOA�\�/]�|X|Z5L}p�.�|>v�H�O��X���	����ş�C��hT�j��0~���m[QG3:�g��k���N�V�wV�H;Q�^�X�ˡ-��O2YM�o"�ꁦ��07����S�B*ji�T%#��(���roDڬ���侫�A����8|qqdv�a����H��%1F�B���J_�Q��L���Ys����T^/��y��-�)�
�qy��2�S�%u�k2J0�����$�pO�6��sd���N��Y�!8hҺJ�����hE/X7���T������D�W.@�B;��&~��/kB$�,ȃ���mN!Cp����bӱw����]�
�L0J�b�uR�+����-�t�����u��"a3&�˝�"�2�1����uUn�1���-�!|U�[(�-�L܃/x���w����?�Yes��
��_�d�q�h�ڳ�q���e͓�<i3r���.��k�;W�_5F�����\�w�^�`�}�qE��,�R-՗����g�ǵ�X��J<%g�+�^�l��oVОx�����N�}����4�h�Z
�D�mo��ֳ��k�0q$厖����䢪D�&|�*=$����$�U[�|����n�Y��nv�i?N,&���R٢-n=Zì'y� ~:���$�ls�n��PA�����@�]�� �~�@xK
��r�6���褴�B�>�Sԍ������W$���$Q�m�O����B��%	��9�T\�3{�5;ē�bj�u�8TR�K���o�a��U��S���G�Ʀ �w�@ހ����c	���o�&��,����ܭE�LI�K}�x�x|����I�OIc�Wʫ�YUޘ]-��M�T-��-�r�Y6�����x}�+��dn�:>eo?� �E�ʸ9��*p����T���PX�����ܣ�=��	�j��l³G��c�uEȪ�|�����}{���o���@o�SiơvFm4k��jO�OO�c^:�D0�e477g�!��q���K)�Ԏm��My��j:��l��h�5��f�k&tN�|Vf�$�V��nǠ��ѓS-�՞[�褣��`_M9{� ���
`l0�f�����d���9>�2��$E^��s,�l1�?B5}UZ�\�^b��>��[����k�;���u�4��3�sϤ���>aau;q6��ck��V�E��W:l�e��X���ly}�T �I���G Ϩ��|�`o��a���W^�q=a1���O����8,�2�7o�X�:��+R[NR�v��ұ��Q{���a�&�Xl
��_&�Y�I���ٙ)a��yi3�`�Tp�ʠI�u���r�ol��(�,\��d���*F��v��d&���a4V�q��EA���A�h�i��ā���
w�������F���D%C�n< ��)���y�\$�P��^X���
8�x���>.{�	��ìS�V6[z\��X.�R��Q����)q�r�놃. 'R���֭�H��K�#���ꂂqC~�D��]��`r�#۱ҍ�Ý��5|����S�e�F%Tg&�$)X�:���fj���M���Ig�8��d��� K,�.uĵ�oU���k]c~������2)�f;بx�;^s3�,,�˴��3ȳ^��`c��qYC ��Q��֋{	8*Nf���wm�.�� ӑ�Z�hw��`K�/�37��d�"g{1+����ͪ�j�p����g�<C���}��\ER��5�+l�;�z��0�׈3�e�\�8UK Cs�Tj��S����-I3W�N��o޳6Lw߭��n��ݕa��_�6)���;g���b���)���l�B��\�B��_~���v�b
6��{��jI��`��r��$��@6Lf×G�Sؓ�3�ձ�v��qyvR�V
�*�ļʹl2}a�/C:gTB�ʳ���TM�<�z9R5�إh)��FM������@#%&�W?)��T��J@�&��x��6���k�7��`���t?*����N���� �,$-Rӕ�x�Y�7擔6b'	QQ���q��ޤ[��+J�f�>�LMJ��7�������+G	
 n�YEg8���j4D$�ҪǼC²�3A͆���uX��1�,�V`g��Sg��P�|	�E A@�[�5���a$�����Sžj�7r��[H�$�v����
XE���m7w��� ;N�֕xq"!��܆�z����Ϫ5#y�����4���� �G����2�ֺ���JO�j��"L����|���½��ŝջ#.E
����0 ���\��j�>4�@*��y��g:>'���d�W��m{�w�s�ԛl|���H�u��<�9`ᴕ�ZӾ�HT����aJ��vNbib��(� 	"�߄s�l��� �c�Y���闳�L�;�(��f�(T*l8q�x��g`���LT��\�!�׻��+((��D�A��^�����))��-��о��7��E�:7�;���P�7d7�ش��������^m`M��L.��`
�UGc�.?[��HU�'|���J�7^����C

H�[�Ei�
c�t�Q�*��(*�嫼������f\�����&B,փ?�7<rr���|��4�̶s�yI��0'���0!q��[˱Y%q�wW"�բ�a�!�BL.��^R�!��x����7
l_I�)7ۓ ��{,�ux��Uk�1��t�x3*']G�P���S%"}gy06�
�
p���<����FO�.G��������>4���I�w���ci/�E����07�p<��[�I���=1� Z^n��Vs���+�,7L~<�k�9�<���E�"�d43�4���q���W�Q�^����޵;2�ٰ%ʱLv
d����DC���s LC���
5�p̷���k�y>�{�n.ݯ��k�<�y}3�|����g���t��R����҅������MVɂ>��2��EAuV��}�.Q�2��\}�@��b�$ ao�e�@b1�o�G�F�����2s�=�qMB@�⫹<%�}{����]�^�D����[�@� %�4B��C;XH��o�WK��vE�n�"���dŤo�G�؍�鏗��d�c�Z�jHٱ@��'���GgRWt�W���=��O���9D(i��ٰ�J��h��w25�){���KFdu����_���	���Z:u�e�3�����ܒj�lT�7)D٨FvZ�[�x3�W�c�Dh�R��x|��r}����;���^�RI�jZ��������~B���v���Y�����&��{7�c�T�����|����w~C�5yR��T��M�]�\O�+�S����������žTY���˙ ��6������$0\8�#�t�y~��㞠�3�f�NDw	�t<���Tc�:B3�2�on!�}���H-�9>�� �-4S���X9	9�I��0ޜmW��J''�ZS��,��|��q�!��� ���ޘuP&����I�5����Xs5O��~�nd*c����8e��S���w�ư�k~�n!`ܳk��v��<�#�4�v}"?[.sɏ*!x�<hi��`�H M�(ߘk")T)�o�/}����&ù�����zU���^��o�Y��#�F�F��O2��=`���*�_ʛ��]�<&'��;j��. jS��C�tz�����t�h�6�a��/k�t�,�U�Ӹ�D����$]\�N��m���oV�眒�ⰰ���AFi��JCkP�f�7 ߞ}q1�� �T�յ޼�`>���|o����`Ô��$[����8ظw��1��
ߣ�&�/k�_�Ҕ�C
��Ў�R[k)�[�	�Ր�I����X�И�6���<�}�w,#�;�q��z���T����vG�
�T"���D�����6��j��<�"���hP����k����^=���;XS�0�o3�Ϸgҭ}��NA�P�{��r��������?Ȁn���5���PV���x$YbO�����c����
��ޤW�̬ 2��u+'7�%�
�S~��/����71Q Ji��Q�g�}�?X9�
v�=x��v�I�Y1lz���ai#�3\�V椅"��i�Bخz�(�)+H���$[tm�u����.}��h��7xO:r��e�m���rNK���SJ�eED��-�YkDB'��0�����v��z^�o+))Vxd�	 }��u����*�݇6[]]E�;^@�Y����1�^&��D 4�1�UC�t�[�SԬ�~շ������&�rO8�Y��?���צ��ԡ��,|{�O���?4^U�����fQ��e=�X���,w��:�zpU�����#�_m���N(d��Q�*l�)��L>�w7*$$��P�uf�d,eä�5G��qq�) k����=`s\���x	>ܿ2\��]��h�s��|��F�t"_+3 y���*���c.�	�V���u$��&zYjǣy�=�г ��|^��ǝT"�{�-\�b[����H$ *�777��qڮD�W���'�u6���>�լ96e�6$_h����߿����Lk�dd�*c@��X�y�nݺ�8�MD^QQ�^��h,iﬦ��N���,�G��v��8�AB�RJ��Ʌc�Ō��<�T�}X]��u��jfHDkC6���hU[�+K7@�@��i��dd��6sݿ�^(---d!��dW�[�4[�Ϯ���'9c�ӓC@.���˫������{�,'���fA�k�N�a������Հ�)�n����{L���`'9s��ԏώ�;� ǯ�[�E3�s8o�ˤ�_��r�9�Rб���!�kT<x�d�_�-�	v?(��$B���c�,���`[Yx�i�s-�>��H��B�c��'�<g��,`pD����$5ł��'Ǉ˭��B'�;o��m��� /1����e�05u�6�U\~|�@���K�U�S��a>����s��"-բ�Vl�Řu;�m����6�y�j�ބS�ˡm*�t����rVf��Xvvv+��P� <C2tr�#�J�� 8S ��vNN�a�=}��ꨒx���bD1�G�b8-SFFF��	8'��m38���5�M\�u�73
G�å��SR��<161a�����Ύ����?��Ossr`�v4Am:�>  �u�L<i7|+��mo��.�]"�~e�J�;=';�Eĕ���4�"�Ѱ��.}��Ԥ*L�S���S߻��K�r!��!� �R�.���L����1�F!����צ�� K�Ml*12|�E8����\2�Z�n��U����R�����k��E!�������>@��� �gȍVGʅK���v�� ��B}�gJF0��T�I��8l5��/(��ʋM�N<�E��/�!d��㫝�YN)����C�����G�������#����|H�EP�n��O�t� �y�r���w���G������~�ip����)cO_�7a��p@�G�n��H�zhՖw�W�dt��1�m�}*�z-�л�oٮ�0��W��R�}뢼�-:c`�4HI�߹ ݏ�S�X�}� �X�~w �LIX||�l��.�3�-�[2�тg�d�ƕ���v���Y?6�B�da�!��tTk �e��^�[e����}`�*�����<K��kԩ����n����j*�8�zxu
�1����w���\�O3T>|@S�D/	���b��v{�J���_<Z��ݻ���SIu=F=����<o`L�����h�7<f�û�s}�����ܫ������d�M�/p��ڱ�����������A|D�T��:�(��KE%����c��p�l�zhR��{�
�n@o�@_�����-e�
��5;����H�8Ȓ�A|��%_����.�+4/���{�V�����5��&�;�Ik_�K�޺����A����~��eٴ��x4�t�k�b#Bm�������f��,�?g�l��꠶��,.�<�%�6��_t���o���$*+�/�"W@8���XG!Wт?Tf'i 5	+�p��,Л��Zz�� �#�,7e���'1�/	�K4���\���/�%^� J����4-~
�a��$�J]��K���)�/B�j���a�2Ia��J3]l���v|���E��n	���
�65gT��R�n���YA�X�&gk[�aU��v�lBXX��S��#�޻�8ᴎ����o^���g�DoU	D]&"C+���+�X�Q쪲|X:6���͘@t�V�4n֚��%ͅh�6�t�m���"͐��sa�tc��5�,��|~�Z$g���9�`���]j���5l�+̂��u�`�2�[�ט������8.�Yl��t�)��w�1��j^�b_�ÂJ.<L3�0���Q�������D�;H�V�(�=3�k���4���g�@�Ʈ}r�p���7��:`;eն$���B�S�!����n��!��a�X1r	#��v�4"�?�&s�4�j�꠆&������-�?���_6,gV(Wm�R+q�S')���+'r�L���� �*�[��%yYV��i�J�o��@�z.�w�9?�p��_UG��Wp�;P:�M!�)b�J#��~-�4;�-����*�/~:��k�e���*Jp3|%��sf������V��g!��	���F�QI'�-��F�ᕓ�j 
fP�?s)��aq�F��_Z�Ӎ�T����'<t��u�+jʖ?�ֺ�[]󕎐��<0��<�歾�X��i��\�f��3�xO�ioQfߞ��0���	9���#9�o��e�u�Kw��)6_��UسY��u��d[	�� ��j�H�ؽ��a�h�C��z�Mc��0��=��.N�gV��* �@��kT�3��=0.J)y{��'��F�r�6VUM-`��e�fi�������*1��4��G�1r�Hǲj0[����"t�T��۔�𹂎��r�Ɂ������p���_�X��y&g�0"����C��c?#9��]\�1.���>-x�59���l���ݒ�+�#Y���7g�v�f7�%D���|9��&�ͳ�=W��ښr;��X3f%:;[ҥz���ڗ ���H}�Rk�E��r�����98��Vm�+F����ҁ�(]��R�W��R�(���E�6azc[�&�=����@v{Ip-��!��!@N�h$�UW^��oJ�V�6�,g���y4&�����>�	#9C�"��b�D���=B���(��&�3�����ǝh������m�ćP0�[,�s�4N��|>Ȍ����HwY ��<ŕf*��r]�I�4�ˡ�x�a�~�	F����r>������"Ξ�ѵ�e�F�Zn��D�;0m-|���eg&�����A�kv�����1Wi/�������}�^�*K�Q�U��H�a��C�%5�Jok)��ֵ�;�=O�:8?�1��26�\n��3FRJD%�����B(�FW=�j[��B�� )ɨ`dd�w���\>XH� tٲ�݀O)�^4����(ۓ�^��8��<�=�<Ӹ,#W�s���A�8Z@�ى�� �Uת�v������3��'<��'�����TUc�N� pPH�"5]ă�~�����Z��0�x��F�����Vs9yeZ��#=9�y[dz�s�vHZ�7b@,�0�Zo�GF��U�o�Ef���>`ym+��[&��B'IVLd�Y��g���L�9��u<G� V(c�-��U"8'�E����I�/�����&������,_�=R�!S���@�ՅG����9	�䨖gת���eW����4ߖz���X�
%0�o¤�
�6&&�F�T۶�ɵ�?+��GL�a��e���O}� ��L��ϟ?�iy����������a���j��:S�rT�k_�ٿ�X?TMp�"&$�O޺��@Z�I�B��u÷W}�m;3J�� �Tb��qr�o�o���C%o�/�#�!�T�vt�,��	����[ 2BR��w�� w�!�S���=��-��x�MO!���*�A-��"��X�����g�r����KbqHa�ƚN��Af���*�Fdy�Ob�����͹�p ��W5B¢p11ج�%���zݽ�(����M���i�� ��EdL[���>�LB�9���Q21tɣ������?�)�����"+#�C���#[B���J���$+�d�B��Ce{��{��p���������Ox�_㺞����%L2{���Q+�/oe{������g��%:�I��>_�/�2-/.�J��D��}A�P�@��-�
DB�9/N�n.�&jpW��A�����z�B��5��@dٴ��.g&����YW���O���:�k2Mۣb�k�O�]&?C���|⽤�m>+$����s�F��"����S*-��>+�+qH�;pܠX��G�=a�`��H��}ҍ�"z�Ϗ�������|�d�����3ƚ��΂i\�����������	��w�*�����"�O}��ج|���Vg��5r������T��;�����ȉk�`�3]�~hbz�wu{g~=ñ��JN��N�Z�!����o����� ��������=�!�-�z��x71����aULX��,�ӗY��Z:�im�n'��Y ���"`�4;;�M���b�kHYYY^��#����,Gj2Ra�p{o��:���jl�(�/��Gq�'�}�l=R�a>��ʌ���)�8���o`� ��x>��3�juk?<��<#��8�a�50{����vk�bY4�@a���`P��~_�*;�[`W�]nCxs;��X�x�va_�c>ctz@�-����:[�w�0�2��00��H*ݲ���bJ&�&�*S�V�4 V~Na�o����\� C���\��/�����a�2�ĕ��� �*�7GQ�J�"�:��������E�1�ʅ�u��W�[t3欏dv���j�х��=Jh[����վ3���p
�E+x�<װ�@����&�,�>�����<�*�9`n��� ��-AA-A�s8�U�ik���%Fz��q�b���[;���J0�����7�p���������4`�tB ��Q�A���@���Y�O7�/߇6� י���=�I��f�ǼD<lſ<}�8��tU`Xϡ��3��UJJ�3�ev�qx}�y��~@�"�[C�WW���� ev�4=p�Xe�N�bh�~b��G�s:z�B�,S��b�9m�Tm�r-���z�%�x�=F;E@��O�zb��V�+����s ���ϣ�P`$���\LFJ?�H<��`�ң QXBs�Lz�E����}��!����q���ϝ�����,�l`�qz�q=���qH�Bp�;W͒��F���t^t�-?Yo��0��XD�^�N�,�f#C}[�L���ɭ0�o�V~��<�<��a�y�� vWvN�c�מ�C�Ik&ֈ���`�VIÜ?O ���l����{���D!��P�)�=��	�v�SC֚(�b���ᮉ�9�5����&��Mb[��������P�̂�Lz��AM�B&��/87!>�=�� 9�y�5;��|o]��7��5���"Y9_:T�8!���LA��� E�(� ���C0�����	�i�Q<�>qY|������V�����$�2��u�q�@$֦��	t�-g+�_%�h}A���̑�8n^����d��硸J�r,D���P��ù���fg��?th�����KM���Do؋�)�0��6Ő���5��y�B���~-r����:�Ϋ�N�6���T$���R)G��v���d���S5BW�q�1'�ө�����w+��,�wi�î����'�b�+��lzlF�$M.��K����e�����_g}���Fύ�B)��
!��Y�<�ߒ��
?؅o���A	�/���l�|�[�"��W*Q���
/d2��;1U��Yέ�]�=M�f����#�Qz&"��[��17$BZ�ʲ���r��BG6è{����t����"ց��xڄ����՟Յ�
��^�\���g3��-�i)��"��.N�!�g�9������vW�Ӕ"���_� l��������XJh�4��-s\�K��z����4M��Ϲ]����Jo��*�ś�
(2R�����<�%
#d����]����뼪)�oF���+���zR���OK�CI�����j\��~h�p"I�^��jio[���sM댋l�k<����e�=˸����鄪�:;�No�W���s��m�#ƃ��Yj3J�)�����dHl��z�u�Z�3h8�7 ����8��=L��
	��Z?��5�鱈/U�w~cK�R%%f��8u%w���:�.7�����UN�z�+�r����-6�Sn���0�R:{CJ���1�p���2�z�����I=R�H����Gr+�S��aO'w����ON�cS�΀�o���N�l�_��t��e�~��+�&ë��:�L��>Y�)��/�|�d}�M9�D>X���M\#F�i�hY齡,Ów��ev��]4��'oEۖA�{��cA�VV|�ǩ[��g{_GI���*v����Y��M�1W�[���Υ3�=���2�f"Vx՜��\���� C�1xsd$����������M�[2&Bme���P�ld� )�r���C��s�o~@�@j}�����q 1�Ǽ��0�_�r�(ի;�0��g��N+��$B���L��|j �T�˿Q�ѺҀ���S�{�lٟ��+���jc��"9��'�H���^�a8�M����ٹ9�Y1��߽�S3�̌��5Uݻ
*rCW�ߚK������?L���x?j"�!sG�c�uGw�2����w�e�V�b��|fJq$RǏ�˘�<b.��l�\�,/��_g��S��zU)�������Z�ܷgY�+�x��G@C���I;�$�3Y�Z��ڨ�a�5B���D�'Ӿ�癶ju<û�J�:h����`�*7�\�~ޱ��������PV[�w�'Y�w�v���J���;���g _�<�3�8zp����mKz��/��ٝf>�,~�ok�i�R�{dᖓ.6*�G�oEp���cޝ�)	Ģ���T���TB�L_΅�_־�u�(I����-�^�+qn�$�hVi���cd�7R�#��[���'=��ai�b�%�U��~����(�3��hͳ�ҔO��`)"�Σ(3О�S�WįH@��Cȝ��jdl[܌�������]�3�������M<�~�b��OT��w0�\�B6"v��T'�IOV�Mm~/u�a������m"=���Ԩ�Q���d�D�R@~�ku�:��?�xN(ׁ�,��ғ|v�m~�F�5`O*��uKƤ ��l(x�P�V]W7Cg�˃�ub.] ���"w�y�Z���fTAEҮ�ˁڪh(��h*���e��S[M��T��l�i�u�\T���5-.K�-�:36������8	�t���w@�� �}JW��9��SV�r&�a��ye���n�WIz���v��S|�N3 c
G/<uSz��B�ҁ(�|��IA��ʚM��a���z7M��#;-���V�r�[�D�����A{Oׅ�,��j��h��Vn�t*q�ׁ��cn�KٺA(Z_�`;/�~^�����������W�b�~��ZjwO��W�+�bq�B��L����&V�Va�Ǔ�We�J���3~8�Q?��x	ߵ�����7>(qj[���d�,v_~9}�τ]~�D�0�v�ѕP�n�l����/�G�ϖ^�r�aC�#�:��ٞ�E��?bDu��l8:���$�f��-!�s�,�����aBtt;8;;�y�(�n���$9����������k��u���!wk��4w�$ux�R�0��C��4K��%��c�%���Ș,���/D�|����dO�#��y��+H2�W,�e��B�W�36����Q��F ���[����b̮�sC ���мN���e"r��Q���WT��ԙ�z3�����L?��ˬ��_���1-�Ztʺ1�f�5�����GL���#���<6���C<N�]j�P��)�G3ї��2�� ˬd&����zL��NOtm����;�;�X�}�g���j�E�ZTO��ﲔsB��ܔ����?�B�8��#�h:Pq����b	햳��ۜ-���m�huo�v�ie�wX(*y�e&`G��w��&Rr,�0R��`�����L��:��v��s�@��k 8�:88(?;I����f���u�����  9�n�&�1�d�����^v��D6��M}�%�&;G��)[��2�z��z-S*�	n^u�RȎ��"��@22���	� ���)'���Lh� 11��45� �j�,�93?ϟx��o-`�1`�~}L�FJF���DL��Y�%=�ff[���-���F����N����r�6�yxW<,�z�J�:��T:|�V�M wblX���\K ��T|��p�4J]	`���7����݆�����DFD ���ӯ����W�H�ae �ee^ �\h�km�1�ѕ��/n����K�9x�o��x�%��
�񥮭c�9����Aw�Z�$�N��l~�TQ��Ȕ��@oW�|��/<��a�H÷��%ϊ1U�mjRq�z-THc�{#,f��JJJ<�
Znz���HU8e2<]�C/��͈`��K=O�OzN��R��.����U$0dc=��lN�:��={&?5b?�bt�v���W� �Q;�7�����?�q�_�b�6��@�o��z��Ib�e��U����(��]����
�u�������*�Z:��"q� � �9���TO�8��Y��Xʷ3%N?o�GJ��Dw�n!
P�څ�7@]t��T�(K��ΰ��(yæ^F����?t���}��5{�
=[���\2P,;�v�r���z����N�Y9����ɓ�!�y�ZCKk6�ed�~�1g �e[�m�elY%,������[�;���.4�6:�p��!���w M���=���;4��"o
�s���-'uT��?&q��9(�Z�?�䕏9cR��g�Ie��֚����AZ�{��c�1|�kYl�Y��8|*���D��ї{���y������9�Od�nӼ���dX�����5i`c��&8,�`lS!+�-���b28̼"-�w	�H��o�.j+��`�*('X��L��u�������3���0�@Rf)=�M�����^rQ�9t�[B��X��!r���ϽC�7�31{� ����{�n'�\b���L�y�.�����T�*�f-֟}��'��];b�ya�#�=���yQȚo��y����**)$�O�]�*�펏��%��m�J��ws1�	aY���fE�����h��q�����X��L��.�s
�x�h�(�W��,����~��aǅ�\`����V�9���S� �w!�*霿��p,��JV��O`/���.��O�o�C*�y��w$ͨ�\|5��&��~h�)�Ce�[�c@,�q떲��ّ �t&{{�xl�g��8��͊^� 9��f�x9�y^��4g;�%�% ��S2} OEYݩ�Y�L�g�]Y{��7g�sF;��[Zx1����ފ���gB�gvf�a��V1�����Mp�+6�AU5�/���"�3�fm��(!;��&^�,��Z���f�K�����������A���6�5� jd�z�T��K�d��B��)��!x;��j��.�ٱ��8+��bCy�'�P����ٝ�S�U���aΪ�K�	-��q)KD'/�� �D�� 
��\�g��G����Ml\�)׼���������� .B-@y�A��?�V�.V7F"U�)��F�0F�ʘ��ˈ�Tl'���V���D�,W�T��
�ǀz�H��)�I=�I���.>�'ru.�:�˪��W����r�y#����d���w�B��X���	>?6 ����U���Gd��і���)6�`	+�T�[Ұm���,�n���墓����h�u���Di��}�������E�h���T}����آ=�<i5 �����r�"n 	QF<OD�Xe� q�t���ۡ�^�̀��>��q�����ωS5��ru@Lk
2br_
��q��	hO���0b�I	ߢ�z��U��##�L"��Y�Z�y�ށx���o�{#O��j�1'��p�b4PVY��C g����Eh����wS�R R{8�Y�)����s.�w`S�~��r�l\�I(�uQ�����=��*���S~ĉ�d��]9�},ਗ��|j�?��2oe�y��W2jkG��׿��jI쟋4j��Ѷ�l�f��<�rL�}�c'A��k�*=i���Zg����1�c��Et�B�xGcm�����_�z>�����X��P���;0`!B�؄�VꚚ�p`�}���E��*���*�uB2���Gm<H&��a瘝de{#8*T ���">��zWbs��`�z�JWR���E%Kp�'�{FQ���3�r9���_���)\8 �tr�,�?m�8X�D����-c�Ȝ �F��Rd�4�y3�3J�	��@`ݕoed�1���*�dK~6}�5�Im�>��3�%�����s�F�5q�wh�}����g�<�*++��6m�4�I��ϐaUL��K/����u�iSm�^�NK��Uj���Y�~���pҀ�v�1B�Uu%�v�r}�cH�Q��@�K ����/Nk!ߌ<�nQ�KJ1Y��@g�982a�'B�Tn1&>3~�E�{���V"�jڍ!Z���IO6w���)8$w�)��9e���T�:��	Ł  �wfx��'m��H�x�;ʴ���b�t����)3�[L��b/��,,�<R�����f��`%:��`wB++E�����e����«��x�퉒ף'F�דn��_r��7,;W��R��I���9�p�RK�UU��I*}�+,���3�t�f���J\�o�����}��p�
�a�,��yW�����w�=q�Ny��+�������v^w1�!}b"q�����%Zú.�5�����NCA%6��U�/v��E�����'4����;(ȕb�?�Qc��/_L���V�`D��n�r0�� �����m��,ws,����`��R���ի�����e�U�����y���̠�i�����>���V�r��/:��aVB� r:_(8����8�y`@�BZ֛(��/�m����xxT�o��pLzo�g�����̨F7f�NFX���7�����g��-ʰ9����h�v3?��z���|�`���	ۄ��(�ͬo)�}~��ou�d�	*n���_=�<��1��y3��W�c����@�4J���k�?�㯜�Α���>��6P`Qd9hp��*�A�w&�ܠHb'����RZE��S��j�O�*�����pv��sX�y�8o��Eg5Y,\"��'T\�0_��а�u�$��]3�%�+�g��9@Q�g���A'1��*�X�Y��4[�>��#ȕ(ޚNb��}譌�[�'2Zk�DzzN��Y��MH��?�8���e����M� ��½��It�-@�h�.\����?�k�N�|��QF�_�,����C� �����fx9s�-U*��h�3 �L��3�,ޱ:�cu9\�D~��	����]�z�b�_܈{�ϴU=R	�-�,�Ɛ�W�
�-���UZ�EɛJ�n���SH���P�{ҩ]]\v�'� ���Gu���? k|�e�}.��ا"!dC�(d���|�V?��`L��4=�S�L��z!�b�<�F���0g��'�a���Z>К�\�i{]/�S@�%�@��D�l�v�ۮ��k2\���ˏ9�IД�\���e�N,�����E�!����wXXi��z�0��NS���w[˩H5�\��P����ɒ�4��Fj���(�)`	�хo���7+^)�j�q!�l��#u���T1	�1�{vL������BH�Ӊe���r^�l�%zw�c�)ʈ8����3Կb�5���`g�����c1�Ghr7(8C^���DCQ���h�&RK�o��\.�M�F*��P����q�� �":ь�:{yE�k�R;w��T�BN���|��o�K����w��*�M9=I��P랤�q�e����8Յ���� �'VT�V��|���m���C�$(5WH��:�+6���5����:����7Cq�p�;%5]��eu������a��v^�k��(k�K���0�.:�%.��{�^^��<�?�;�(��z�2�)E�3ݙ�c�o4�bt�'zlL׆G��ʤd��n�h��}��Z�QOgvuY7]�;0��
I,{�l��w�s�0ǻ��6!FmB`p�����*����v� 2�g�p�τ��v>���^4�K~\6��Mf�����3�Cy88h*BR"ZvjPM��&f�������Z��O|�S��P-c��P�>p���r%k���A���	���Aɇ{S+�5��U��`?�l���WR+;���u�w���C��X3{=��5��p�]�����T����[59��W�Adt4Th˗��S�6�����⽿u6q�r��(��ɒx��zF�>C��͇>�~|��Gva��P���pq�]X��QK�%<oؾ�5�d�&��YG�O�ݐ�줺Ȉ�3!D�;����YU��쪻�qI��r��-_rz���n��H[5�\O
=ձ���R,*Q�cM)��-x�5R3A%��r6V7u�hފ�b�b���� ,Tc%O�3�0���=�x���oԅ�y��@�ؓ�fv���^����V��SI�OzP���aH���k�Ū#�&׻�U7��!�w�2�� Z�MI��T�h힎$����NX�+)�9|5�U�[U':6Pk�Խ�Yu�7�;t%��O�kbx> �)��#�����;���{kY���⁉�o��D�A��,V�*��2�ku��%��]�h��mˬ�)�rC3�鼿K�v��)�>�|��׮�����>K���Lo�<{ȪQ�C���2#4�9�ڣV'�A�����ah���ǀ���^ס޻p�B\��bML���1o��-���a�;�;��֗�Dֺ��N�Rw~-"ߒP��<v����h���8�R�r���E�;�N��>��iZ��T��wN?��w���c.���ٌ2+T�ߓ.���X��:�.���J>�9+q��B�p����"0�F�d2�;s�9S�>��.�h7�?�H�$ͮ�p����g.A�x-�Y$���`u��f�F,��XJBM8;��M�s���ֻcM�)�HY����������.T���{vʻ^^U���1g��"j*h�[��h!��U]���;�����������#�����+_cc�*E=`*��c���'ۥQ�T+v�#ʱ�(�E[���<�����S$�>Ć�ͻ��%��}�j�~��%���Ӛ<؜Z@�X�D�n���1���]��\��,�Xhcq�� ���h)��ai##P���no�S-t��qƭ��rx�*��Jm��=�El̆'��J K�7�^��������l�LD���%�Fh�s����lBǻ�6<���������oB�՜��ϕ�]p��u��Iiw���X���=���+�@� q(8�t��̏����U��ij�yR�����\v"������B�+��٩]�
bO~�]-5�W��K��ڬ;��;u�sr6VVH+D� ���~*�����wH�K;Eٲѝ�9�(}^��g	q�:؄RNzc�6� aN���P��@}��>At��!|��.Z��o�}}���B��S��)�>1�2���	]<�tL���V�n�F�������Sח��(7	1�Q]��<�)T����o!��͢�ػ� �U�k_ϸ��9���1so
�CbB$%-x&sb{*5Wgwi�}�������J���!g��y���ꮞ���֝���<F�|?�ɥ1]��Mu�`C�pxv&�E�]rz��tVfRO ��qgWW���`�]r�HubG� �[t����SI��5^����7��u�e]0߸����X����	������BH�d�A�&�'k:v����6��B�-,��P{�32�.\�03;�fe�s��7��Or��H��ܢΞ�,5~����f��H�.��m|f,3P!$>�el��-����Sd�WN�(^@	������$1/ys��������[l�S
�b�f�}��2Y]B�%R���^Cؤ��:f���LJ
B5�u�t�A��C��Dq8j��N��b3�PR�w(�>��u���ԯ�Q��=KD�����<ۄb���obUu��j�.����´ֵh��kGO���',-��z/xGo�F�q�������b�z�f���L��WF҈>����DHrÌ>�n
�\�"Q7����1��>�7la�����d.�a��^��tIH��x�G��V�����eG�?��e����3S2����Md/	nt�E>��|n���?�4w	3�6��F}ԟ�Z�-G*��R�N�����CX�3u�i�`��d��|2Г53ە����JҍL��QUU�B�����KO�n�X\�v83U����ח��6��;�iiD�B:9��	��U<��p����	oJ`;�u�jQ���[���~�mиw�=��Y��)HgR���ֹ0�j�K
N!d�FM�	��_�K�^ M�D�Hf"舢.u�4X�&{.�ѯ�79�i��掿���rc�K<�Pp�:�|�� �ŝ�@{ߏ��5Y�M�kw�AkJy��<���^�����p����|��[Ӧȵ�[� ��v�?��B���4�h*�j�?�,��9������P���e�%T�{}�����GKf����!�Tm[ՙ��m��r`�U�(���4O�J�Q�ۙ�[�C��P�����b���}w��+��<y8����w�⺫9$Jn�篣(���S|����;9_��s�y
U����:���6 =~��^�޾v�S�=M|	�h��*n)�Z��5v9^�ﺙ�K�C\1�>4mţ� G�o����{�X��S�D���m�7t��U:����Qe�L&�/�*��.��>w.} <آ/��v��W�O|�'1<����G��� �����Ҁ�`����&�;�)����ڋ��������h�R=h����Js��JO ���E��e��3F��?��v3��U�����pC��[�*_��D�O�wۉKh�E���"i�_,YCE-��^az�T�h���Q��eT�"��6^@��sor�c��@��'�1��쏇�W.�(��/j�x�$?��}�V��9X�2&����jv�o1ﺑH$�G�S���^Ȣ:Q])��/�a�|�⑈� _��� E���*�i��<���M�+v$N�{u�<Bt��48I����n�@;@�I  �E9:E+���,�(_,���5�����HO�����ϓ%^bQ�KK��
���CT���C�{u���m/!�^�R�h Eh��\_�?Y�����s�<G~\��2���-�]��z���)@�Aiii��_C����ō������o��>6�<����8�D7��V"d�.��kc�3(���U������z∫h��[��P��P aL�y�� U�o�tU��˖;Lј{��+,�6�p��6�����������򙁯/ٖ߁����8��^u��?�^���[Z��"���m�{�x�$���p�H��b)��Q��A7`OP��e��d���Q�v��o ���[&��A���+�gQ��y�D�G���
|�(�o�K�NļI]C�bgj�4��ֶv%��:p��x����a���ۭ�v���q�:���'��${,4B�.��?T�ڟ���;���ݟ��[|usf�Rl��";?� �p�^h���V���i�`/Y��호��|�S9�(6��ϝ���*��
ȱ)��`���7�y��������l��b��^��ӯ�g�V
��C�yh[T���\Q{|G�]�<����<���.3Yp�$"�G16t6������Qr"��є[-ŏ�'	�i�q�@M�~��-K_v_��E&<]��6���<�@tdDD��fDDtgfn���صޝ򿔚�@�fs��qs{��[j	\,��ߑ�7+�S8{�>|]�9D���
Sg�X$�e�^
C���=��s2���
���N�bI��:�O����W�� � W��7��{Ac��I]vx��4*���'���Ipk�e?e�\P����JL�E��ܟ��65�B��96 @hv�ڵ�ƹ텤�UwY��� H�̬Z��m��'Ђjl��ӫW�b;ө�C��ml;nu9!>{c3��<�N:�rrP��Y�E�.�'w�Z���A� ���H{>�:���ּ�Yڎ��\��T6(�/֓y\:� ��,ߩ�E/��'��nw�?�vtqq����OV���Sc�����j�3��+}��(�A��"��H�R���Ƃ��0�z�X�+ �wp�0=�_���`� ��E�2����}�o�|�!嚹��BE�P˄y;]��N�>��.	R}�zݾjo]2K�����@�0b����"�6[�!��o)�*e�e��Z��mI�aߋ���n��aw=v))����!E@]�s4�z��}1	��ceS�8�K�R콿sL;{�ꍚ��Z;�S��M���۝U>��(N�մ��0D�%|���ahz������Fɇ�\&##өr͓��`~I.�z7tR��{�m�TK��tL��s�/�[PP�b*	Y�9"jv��xP��]��T��L`�T�r�y��9B�*�<R���g��@w^�bB{��SX�|��U%"��:�a��ں��q�5�O(� ��t+��]�wsg�(�7����E�b��'^�1 ���`��0+�+Deq̰`vd�D,?s$%v1`�C]�P3��`���躛+;�
Z��m�]�� ��.]5�X$v3x
�f\)H_�yU�,ɋ��o������2��f���hp,eT�xVb�^>ߡ�����D�7;T���G��s�.�"L�����_�I^"��@w�@���R(���O�c��hm}Ü��2�X������^dԏ�(�Ϊ����D�R��G�n~����YH]���Wd�c�F�!=&���r٨�n���L��$�E:�!_6�'��qOp��ODT���p��u����KLO:_g�"4>}}}���_i��9�`V��? � m��.~�F�P��v���h�?�����!f6ڠ��P=s6�u�eg�H�K���}8`]j�%i����aI�.<��$Յ��Er�&l� ���e���W咥jl��F[5\A�4m6�X\Ϧ��=���S�I����l���<ݲ�*�]����S��dg�P�U@o��F���x�NbF�G;݇�dӝ�l�0�Zlʸ0�XK��T�G����JIF�� �}���n�@����0�0�hɒ�eJ$af�����E�"���;��R��b��a[���,���[F�U ��Ӓ��[N�D�g���w$�&�w����~z��m��0]\��Cx�^���!`��Ȫ�R�Q��P��xC?�I{,�(������%�F�4���"P���Y�(J��������] d�\���mFkk���g�s����e�`<�#C��u���|a�$j`��I�;mU��	���%?��i�qý�B2�������>���{>�j�+;�v6'ͬ�̬¯aj��K�{�C�����G�z��9c�sz��tR$�Ɣ����ܦzVZL��,Ӧ�Z�g���&ɠ��'������N����Nv�#S�.�ZP�����2�������j��Uk�N�P�D�L�BX߱���ή�}�9Z�C|��p�o��T��m���h�2v:#�b�zM:�
��*�kS_nn��ϕ����|��I�?z�^��iw~s܍��]��zz�6F$�^�W���������;�%y��*��U�Jm�V�Ӈ���M�W-���(��/����<?�ǳ�O?��Gw�QM�M�e�OP�F�s�q��%Jҗ���]\0r�;aؓNf|�!�AAA�ۓ�%ƍ���ŝ.Uh(��1`6�@���ٲ�}:�6�1�%����n�F�7���Jɪ<�bM� �������^;͂��m٣�v�`+�I�4��/�}O�6���n��i����%�̴�{[g���j�����w�M�Ug7m����
���Y���7�ܺ7���+�7��7�ݒ��I
�~k���Io9����\����X�)"5`��0���]�]C�7�N�ul�肐ڔ�'&���
	I3a������R ���Ɏx�*��9�W�И����'��/&m�P����:iMp]�����4j�Qt_�Z��9�
��3Ԅ�a��S\&I�o�Sۡ˹А8�Y)y�zh���<��f3�ÇϽ(C�(��e�1a+�o[5/�����1�	JPpa�0�����D�<�9��D�R���1�]�q��A�V���s��,�\�$S�<=noTt-��/��[��3��B��d���s[5�"#�o����)L׽�2D�ա#�|�S
�-�R��#k�(�!�N����gTxyUq��9���;�oO{ҭ��$A���d��0��}vYM#�+�ڽ�{muw��ʭ޾~�켼;6��sH$���y_A����ଜ��w56C�.}j��Z�5ka �.	X�,�a�.P��6��Y;:_���ŭ��-+�J�g���J�ī�f��ҁ�Aے�B�3�vRCKW�
��-���4␰��3tʮє�dJP^}�>n��`����_1}�+��
e�(�M۩l~|����u�5j7�p�,tL�%�9,�	���⽖Z9�_�$%5����ɹg�n�*�g� /���w�JcK������<�����CZ��[��b�>N M��x�nܹ8+���/v��ʫ���F,�^�� ��cϜ��*�A['S��֚v��|�� T���?��9Tf��\ǹ�~F==}���*�.�8@L�ڙ��2�]��˚3%b}տj9Y�_���%��y�hO�4AG��=4��ϭ�,�?������~�5�`��q�F������c�`�}�:��s�{"�k����xl�^z��2��!z��zP�f����Ay�>alY�<ٕ�]7B�r������CϵCP�~Q��Ss"�;& z����O��\K��M�\-nF�v�6��J]έi�A!u�����F�UyYB�1�Y��.�����P8:�`�G�}`�	�f/��_i[t��s�ٴ[>Y���	�� ��uɒ�����rPx�R1dh�h���婏��ξ�4���}%�6�Y��{���gfg�W��~��6M����#/��\l�U
�T��n?�w�ۓ��o����&���t��p3��k�/h�y M���������%�c3g��`jǠ��u��C����-����Bwj8>1��v1Z�^zpX1^1�.�'CPfq&_��=��3�5~��~��b�WJ&��<ֿۓ��Z�4�����n��GA���Ÿc/��\�ը)�N��~�l�3����-J�M#����Sn*���6�o/N�`��2Uy��P�bb(J�zSQ�2&;[N_�{i�}���i�Q�kw��>��==3�O�2U&��>�>��' ���%�[�j;3Zu����wԩ�˯7-�:�a>���%��2�z4؆s���������?s(������H��A����ý26vg-L�_�����������q�5�0,h3�����iY����?�gZ�%_�.����R�[a�&]�@��3�>s�ʤ���ͤ��*�?|#���ڼ�#7�]N:�Xk��11��$}��t+��TZ��g&o�{�e:r]�;a��]���� )�"�v�?��^O�{�x䢯�Wr-ᘤ�S^�M:�l�ӊ{��<?�0xb��f�ǥ}�L��K{�+"��ν�y�m P[��6�h�A}԰�&��0�/y>84�ު�z�j�#����-6�+Wh%[�.��?+�j�z�.^h[��6�'ok���z��-�*��%?C�<���XS�\]_�S����ש�;D��<޸���<���C@Ƈ^ر����>�*�.&[W�{�E�oy��W�vT�_9󸿓hFӈ{+ii�y(�r<$L|�r�(-�������0Z��9>�6���ћ�#��]ö�]"֤�ڂB��}��Mڣ�K[�
�^{��9Co8�2�:k>���r���=��wf��ݫ9�5��}����*�����OB813��b����dʋ�2hƓp�����װ����@���$���@ww��{LD�x�1#��]J"vix37)����s���P�N��03��;&D{>��r��If���`���,��6��󔠹cW�Swݪ�%�����/#��cC�{l#s'�?{ !-.��'��y��g����v��]:vt�*r��d���S�����仉h6�J�Hb��$:et>����ȘH~��x@������u���RbJ:z�kaD�EJ;�n��LU6�}#�[�eͅV߻��#)���MT��%����k�C�q�0[�l�lrgr�X)Rd�����OfnL�C�Ю����'�V�X���Hf~�+5����ݿR�6��plog_����vxp�؉㚩�_f���#UA'�8�+Q+��L�+8����ֻ�͕�|��t��s��j7ۆ�eWKkY�^�Go�%�U�,�Ƨ��E�_QN՜$H:1��_/���'CB�'�8!���b��]����Ȩ�'�/�Gk�$��w_Oo|\�V{�m������Ì�?�f!��U�f�U��R���p0��KZ*��üu��%'n��u@���9UB�2��c�-��A�Ж�]u5�C٣[k+�Q��%��*:S�3^�v��I3ݩ~�?mV*�*��_v��/_���2�^su�������+g�/�
q�b���J��|�j���:l��X��4t�WmJM�K�Q`www.�p2>��0���u���jd�Aى�����Z�ɦz��M��`(��n8T�^����p�XDf�:Y5¹�0�TP$�D�y�{���ܪ�1p�-��,}_�>���L��_���	�
6&���������@T�1ol	
�P(��U��EW�n*;���l��8������5�t�6w4�:T���!���ަ�%~p��Ю�Ҏ�-i\V�e�3�������\O���'�ő�D�Njj��X�� ����\�_=�5aD����#�b�<]t-��?Qi[O@#߭�2.�缮�
�.o���<��SN7a�X���dI��D������B�(X����fՒw"����ɠj�<��;�����ӳ�]���4fz���C��Y��������t9;����W�Ӟ��=�S�h]t�Xo����m���'yJo�v�]�S^x������\j�zp[|Ջ^G�����nv�ޗ�� yN*]�T��<���C���򊉄�}��	���YN`[�}ZU�6�B���QWos7�y�xd�(z�y!��=�o���
n4.�*�I�{�2�g	��}L2�a��jJe�p���y�~2�q���.��q`H���ԝ�C���'�v�f��<i��N��ޮb$����k��w��(k̯�I���#;�C��o��yL%B���oN,)�k�d��k͊�����agƤt�C�}AI���Y0g���������l�Χng����A�T���a��o�M��XS�^���+'1¬��L����y,��}�a�i`����ca͎[�=�t��s6�4�`�6\��R	�6��`��E� �W��^}������z�ݜ��Gl2J��=�J�ʯ��|��)�W��}^�?H�X����M ������r�qs@o�ۍ�Gg�!m�Q6e"�xcU��z�\O׾�u�)뗽���u����f��8*IL*���ۆ,��kDV�}9=7<=ʸ���>��Fte0�`���Ƹ�6=�ホY@��G��'?��ﭼ-�eV���r�a��P6�v�d�;?�?3֔A#�\�gJS����y-0�]�+�C���?y���yI������|Ծ���;a�s�����i��ժW_Reb��s&�{��M�|T����k�vP8�9��]�xR�4N��x���R�'�0��6sa�� �I$3Y��fC��8��4@O�SO����~siD�ˏe��{����/"VYQ�[J�|���:Rk-6~�G+!�I�s���#4�H�R�K4����$���_���|�I�-ł�e@@�t�s5�/x�mQ�y&����#�!+�U��iaw[�N$�Q2w�\�ZV��p�1 �ڦ/?j�p��'X"��N���[����>����{�*��}�xDiRB��PA�D�tw7"-� ��{�Hwwl�κA|y�q�:g�1���ϡc��{͹f\�k��֣DE��f�3�eRp��l��nM�OAzx��P_ʓ�+������|���� �E�f�ա{�&5���Q�5p�dP)���ݽ��R���,�*ׁj(�@�}��c�sq.�zx�>f8��8[�ᢾځ��oV�fR=^�C���4�7��B��?�m��V�7Sor -,�*H��	��{���P+*�Q��Z8�_�E�����>+*���H�	�ߦxJ��O�]Y��7� &���{�D2��N��&��;��ٳ�/�"FC����>Ɵ�N�'�$N]u�xZ~�q[ߖ���(mS�ӕ���F��Lh��٠Uwö~����ڒ���V.���?���̹؟�r�� �N��W(����4w�����A�TE#�}�|����qO���n�k(�濂r����$g�K%�����P�[)n�t��8;��!q�3�&�A�j^3������*��˾�݊-bV�I���d��r�(G�q�X��З*m!��J�P���{vP��-�P]��j�d��dH����I#z�P<��[;��J�ޥ�u��j|�y�+\q�Ml�_o�?>�P-��*�ai�8�����="9?@��$�mI���R4!�b�4���VۇV]��{�O/���:f����)����T�d�8��[����*M��O(7���2m��mt9�h�R�D�� 9q
 |>�xd�C<6!Qv#΃J�|�i#Մ}'��k@ۼ������ǰa�|'�*J��L7F��|k���;Ʌ;^4=�蠖��������I�&�����&'Z��ҥ�|)$�z��U~ h�=ܮ\�8�r~s���5ߖ����W�x+]oA��,��.ETs%(��O�9���H�)�
�-�۹%��1%�rBZch_�{͕8�Yˡ���-��3� ��s���� �mo��._�Ů �� ��݅�R�G�����ғR�(D��(z���>���%Q��X&F�8��#�|�� I�����G�}����U���][��R�i7Y4��?�T�%n�s�z`%��_%I����p��6
jm�/�����
�ՙ�mDH*�2�y{R��QP�`��=��(�9+�1��^d��u\s���/p�׫�0�*n�6������C��g�+���й���@d�a��@���:-�>q�~1>O�n�vm�ɚ`��@�:��Tv��7:Q>��&B�~�����S&Ꮋ�1������OC�xr.diՊ�O ҕ�� l���!.��+�|�8xԸ�zl��3���ťϧ"L 'T����̡21c�� �=��0o����[wvϖ`RW:��� �G���4�Eq������K��˨>�)5�����F�n�ҽR53燖����]^���M�w�#����zH�-O>A��m� z<N�T��4�L|�T�]T�)]R��MC����q^^��~8(+�ֹ����u�D�k.�����l�'��>"��@N�o��"�d�-ǖqlW�2�A���n���h�^�!Ʌ݅X%���{1�R������FO�wv_
��5l���o7�]qZ�	�4�s��`o�TI��U��w�|5�*w^>61����>���	���C��^�9��Jw+����d�t�u�"8ˠ\�`��@Vf�Չ��^�"ǽ��w�`�#FFϝt2���K��|���l�r[�Z8��;��ڮ���s���4�0�١��W� daD�W[jU M������:����NB��Zg����k/������'Gpb]����z1�� �����u���=@k<m��kC�d�A#Yv�κ��O��Vsa^�ɒ�����_E�� �㪖�)
�E�\��R��a/`Im�̛T�e-�X�KUrj�G$жg��M<�4�#���Egz�J�KOLL<���*��d����xĭ�80�u��T	��e=�Y�ό�/�"Lr>��%ut����y���yl�w]�ߔ]�K�Qq"�1ҝx��E�={�{Л$��^e��^'ͦ�T��Y#�/���FW�cG�+��]�zI��2�,�@݀D��Kw�w�w�L��<�ЏWo�&��SY�9�d���R�D��Ǡ��q�:�7�������������B:���`���6��Q�`I_٧�7�ˑ9,#Kj=l,[Lj���E�wP.�g�����`�M�N�!��l�xضg2����@�"�g��A�:�"(%M�M+W(���cM�(x�⹇��ꤔ�ƥd<��e��r{ƺ~������s�
j�nv��	ٽ���sƺEF0w���,�W���*l�ل�/h.�����ʎ6[��gC����@ߑ��6�j�U!�`�����ׁw�
y�g�~���'�B���GOL�1<?!�_BVeu�=4��7���ZDA�yD��Ź^����gӮ �޼�js��s��d�ˑ���:w���|ҭ�r���`v�I9�]8���r�FV��������QL�>�P�G�h��,�c�u��{(6K�{/}���O����>]uZV��^,�UQ�}�����5t�1*�(��5q3_V��D.��;��Y6�4�Ԙ�ta?��Xf�:d�W���>�4�|�~C�Fg�3�4��ڼ=S�Ł�4Vץ�Q��:.���z*����!��~���.����}P��t5k��$�
]��3���8_I*�.��"��ѿl�K/F�>ܾ-��9����JwI������oee���DZo~���92�pKū0��ن�v${qc��[>'��nC�@���ݱ��l{�a�k܄�<d�W�r�=�wz�G��8�x9	#�����G�^+)E�2����dE�zd��[	�
4'���W��+�(2�^��>��t���M	�T��n�4:�Դ�ļ�#��O���	w6N�չ��_i��ƋNSo�#z��e:^�g��-ah�_G�=�-wZ�\r���:��S�]!ϊb</r+��Iѱ)��K��h�/�姊w��_��"aru+��Bկ���9�\�ey>3����%��re�.A�蕷-Ж����U��u����0�K��B����W=l/&��yv�u��N��}&�p�٠aw�kB��h:B
�%��Hz�og0�mm+*�>�:jE[��L�&F��Q3<X@��M�Sg�U�n��t�p%:��r��i=ZV��?�=�C���E{�Ɖ:��xQލ[T����5� -�u�'��4��!T
��\�����M8�w��?�1y6���Xn�_0#ͳ�k?P���]��|��DD1���t|�5w���"��_n}r^�G����F���B=��Z�t�4�d�g<�t1�זw`)J��N���MT�ろ����$�Z�u('��A+*���3�~J�:��G��{����*F���0��'>�{�������F��l�ѥ����֫]>D\ }�D���2�F0R��`��E$��̱���ɸ\[b7m����8��.�r�m���\Nt�o�we���P�ؽ1��;��1/糩��r�bw=��ֆ_R�/�o/�*�Ď_��f���=##Y���#�Uf8�5t�:�F�U��]F���˩K4�u�6��Ҁ�j����ȿm5��RC��e)��t�+���	2�!�R��"��s���B��$n#���b:��?�]�}dr~�	�k�p�Z��")�&= �}��cATis�\�6N�p�M�#�Q��-1��1��T��c��D�S9 �~��Z���[n����-�D�t�.�rT�\.��8W�3�?�x���GZOP���=�hn�3�kW&N�Wx�mf��|��̰L��s��,,�V^/�=��%'t��K��`��!C;k��1��T�ݳx�bޮĐ������g���������I����N����Җ��B-���-٬5a7��?WϿ������[$�H��y+=��>4UL*3�[�V��Ͼ����f\+���WX��</(�Xb���	>45R.�-'-/��7�&x�Ԡ�x_��#*/e`�1�\o`���]ά�_K��uqxQZe�&�������S$�f:�֊v{/���#��ʗ�A>�)�"���jŋ��k�s!�B?oYa40z�J�3K���bQ
G �Z�db�c����D�7�Z�}K�X!�	����WAi�f����~����1u�A��t�lJwJ���[�^��z!�z2��F��;q��J}ͦ�-�JV&�����_l�|̀�^��x�P�:�/i�U��Z!�j2��O7?�*$	�-��d��/�抓8�:ԋ	-*������æ���B{=<�Z��rWM�}Y��q�[
& ca�����u��~�c\+Lf�8vb��~_�f����nW�{� xG4%�ٜT`e��/�����,(�7�����@�z8�����yt�r~봹C���o5c
�͝TvmiNM�?�@4����-}{�U+�~7n��%+W�`F���i
G�\h� ���_��B����䟥���=���F}Ez�H﮾���]��d�j�d:���1Y�I���h����ʬ��+���/�\�l5��؝�k�o��knk�Y�O��&���C����{mk����x���r�hn��vQ��Q��������Ğ�A͆����!J�:��%=%�_ȌjZ�%Z�>��hQ��u�����Z�x��:P�����T������J���6���I4�Y�ae��7��7���"�����ԭ�5�:
4y��hWf*���z/�����s.P�˅u�$�DK}����%2Z%�aB���8H�\���M��EɽP�e�4�Ӝ.����[�;�\������]��6$g���X�)�U�S����?J}�9���[����G��֜�h���9]+�ټf�f+��=R��~����[��.J��t�(�΂�]����vL3֛x7K�td��ʨV�Hs����ʧ-��\�<1�v�߲�|�ꂯx�g���*�|�IG��J�;^� ��uP#�K�]�쮔6�;W�F�u�uIE/tz���~�hjhm�u;,�xI*�n���L�|Ht3MC��'ԝ�bb]���)Y'��ģ��Y?��;t�R�I���]�^�
�{�G+ŧum�޿`k2���U��6�_Oߙ�K�I�c���2v��EaJ,���|�8�6�|�+]��+�<zQ�����'"	4/�M�C3+S�O�+�d>Wv��@'q)F��p�l�$jQ|��%��x���;�n�Y��VϨT[��KO�>�+�\1�5co�����>�Z�A;-D]���\�9�&)��5�lP�5̼0���6�&`L~6b���M�Y�ڷ��o�Ǭ��*�����a �ڥ/��F�?.�sm
/
�"PK��ӐeC�N����P�XD>J)�� �HVv(�9x�k��B���[�w�=��ȏ�Z���B5�W^dF��8�����S���~[RekS�yЭ�tL"�-zX{�4{;��,����t�[�pX���Ո�1G�h�:{�o���<I��2��{+z��9J�G�ǼZ>���M�jw�
���O��	�d�ɴر��B%�.�v��:u�\���4��m���w��G���Y�:�?n���_f^�7�MGU����W(�댻�����^1���J�������~LN{:��E���g�� Pnt/ⳇ�`�u�>���[�e��^���ֽ{�V�����������F�QYHȆ����K�T��yC�Q�[hQ'�)�{��)�x�h���{S��T@�R�q�[yB�J�����J��D��4�W/N���k�Vӳ>꾚�)S������:����PKTJ�����Gۡ�Q�n*�;$�+��Oqt�W���:���V��+�j�9n�OLm�������!b���Z+=@�Sl���D �ќ�_O�r�`�b�����3�{l
L���v��E�j����Kȕi����I+��Ϟ��v5���wI\֚��Q�+ӽ`���6�zG���F�㳫����H�3ϋ��G�h�=��G޽�c�7�E�P*<H�A���6�/�;����՗ȝ9���fg����
Pg���&�65���6�t9��y��W}~�?�� ~�{��`�4?�y_
E���4J������Џ�/���Pgs�-��O϶�d��E�s�s,+�u�Ie�����~cR�N�1��!yx�1�a>�?v��>�CR��D_�=!xQfd�oG�2���2���Z�A�������c�D�櫚�]Wq�	��xSI�k.�c��)����b6�v%?#
f�7�#�2e�k`n�/�5��2�_KG��";P�)�עB<X)r5�,��9ʘ�_�,^�Ę�#Mi�G�r�����:���}E?�1��G��%:�c]Yo]��5S�89Mb@ܬ�?S.���_d�^�����b���P���9/����uТyJ��0�8�h0f���F@����n+,�NQ��cT����?	_l1~4��Aρ&۞��gI��p��c�16wi���n���\��#���5VX��9{�d����-�P�,�]]^�$�T�T�`z��Ov�CD ��3�՜t�\����] ����5�E�t��ѿ�<�S��*��ʿ�a��A��y�'���5k(5הvuTй]$J�V$�j�{Ǽ�n�hnHԘ{�p�]S�)f���elq���_f��w�hk9���1��6Q�����gM�E�8�m���an����b����w�Jnהܖl=�����Dk.d6�;7�M��V��-c"�2ܺ4�v>=C��m���B/�6������u��mّ���s��LS�T��㱊�p����G!��B�����E�HeI�'.s!Y��߹��&?	�愈�+w��%_o��ů��b�/�Ɂ��GY����5f2o���L�9�M�a7��,��w�F�W�ȏ����:�ws��>g���Oyʢ⳼�&�o�����VU��ֲy6�s�_']r�[L��.l&ˌN��]�y�͡��p��	в2\�e�������O^�܅d[n���.��XI�J�>�noP�W:�F���8v�0eT8Z�L��&�|��f��Q�w}���?�\�Յ"#������:���<㿘���5`�_�V$Q��a}��N~�x�u���%0!�5��ȳ�;n^�d��GH.��?R�&�w'�1��^��U;�يDWP�&3Q�~'����,��O�I�R����J�ճϥ����>�ndxu;26e��)]l'3�q�������*��a ����X�s�\���l�U����i��\�>y}�Q�u�[<}�)[r!Z���2�gv���Ꮎ{�CKp̩a����g���-��Z�X/�Q��ǵ�_�&n��6.8d=)g�p��/F���9�8��b������|��,!|M���)hY�����x��<�u�	��z���gA�X��R|/�Bwd/�$׮p(b��{��㋥N��lY<��ao��N��{-���;��v��q�D��x�f��"{x��-���qՃOvz殺��p�1PD�}��g��ʣ�lo\�����]����8��TD����]��'�J_���H��H��Ϧ�Zs�����-�+XF�+C�e��{��̥<6��=���o/�����%��t �����	�#���OU~���@EA�*3�J�ǃ(&���rK=I�K�'msGGW��|����O��p�K�<�n �^&q��c.�8DN��|�r�o����R��pq��x�>:p��N|��H��t\�>�����i#�?��x�"��n ��!J:���˺^�N?�P�2:������1L]�(�q[��Ӗ�o�\���ϡ?d��e:t�%"��2#�f�U�|_7�?Yu�5r�c�����H��9vKr���^��AYxV�0]@��NM-w�^��nUݴ�f��YW��'���q�����+st��p�����{4sn�к�&A]q�J�<�R�B���ZC5���^����M�;Iנ�Y��Ĳ�O��7�5B���r̠���b����� � ���fg�J5q���Q���Ox�,h�� ��jq�%��;Ʀ�$^�8�1\�C�h<����_���f�bJ�6)������g�X[M�l|:t^��v~��w��%'ǹ�2:<�N�q��֯�&_�}Ǹ�_��b/�\��җE_+��6m���?Q�_�[��2P3{�J#<�o��m���5���W3��I^�#}��p�i&K�U�㏶�����s�$����5CG���*�l��r�a;��*�� Ԑ�:�)w��S�&:٠��!�g��lH�^w��m�rF�v�Pٟ���!}�H��*�S�8F�=����˿�9�Y&�:"�^�����{��p��p͵��:�I����7X]?�
G�Yu�Z��$ߔm&�Q��A*q��A�t��4�g�K�k�ی�S��-d0(j�+����//�T��J�F�nR h�(����&�@ި��Mb>#T{o�2K��6�1~�w22s��K���2 ���_��})p��ŭ+��&{�ĪݍWm�Z�,'�a*FC��F�����蛕m��t?���F���v���x������-wǅ]W��hu�u?��.�����G.c>��mC�`��|����D�bǌ��ZZ���<q�|���<�B����O��WH�d��Y�HA��2e풊0Q�j튷w4e�l@��շ�#�+u�k�z[����tkSP�	4g0v�o3ߩ8����M�=�Op�~D�
�ct�)��1�ISOG�8l�ՂS��i5A"_\���@�Jo�2��( u��}�~P���M���g"'���&���OƢ!U)�ChWԾ�}��owq�ߏ����?$
B����A[�!_�؎:�c�J�����$u��������y
'q\4lw&z��bR}/^��E���2�馅�Э����O{!l�<c�����Rs����1�����f���9#GU�)������{c#|�g�"w: �|���m������zL[G�KI<��:F)�3���?2Tc�T��Y�f^��x\��$|k��Ỗ�>I �p2
|�v��	cg�cy�sP��;q�;��~S�o,E����a��NN>DL�"t��W�x��*܈�q�~t|�m�6�����.�A\6�M�6���.��ŇD���������%;���YHn\��Ҁ�,ϑݝ!�� �Pi�$���ѽa#�zL��YvÇk���-���0���~A��>i�-S�V���jP��ȓG�c$a#[���1)�5�گ�?i���.-e�~;n[1?M�����ƌ�0�Å��{�wFg����H�x� ]�X�>f&TW�UjSm`ypT�?zͲ�oӶ�J�7��K��Cou������y��3wT���'�&G��Vq���𴟮.2��V��x�����$���W3�w�4�@L<W�b;��~�mD���DJ����]!I����`��|�M�F}�����,�����ʠŢ�[�Ю,�̀'J<A�|��%
��I��'hǉ���W��D:|`ǵ�+v���|�_��/*N��5�'�	�?|�K-��?���{{h ���D4y��������9�y�Q�걀��=�X�M.'G��j���#��4K���|L����p�rxr����145-� ��V�;��JV7���%�|�"&~zե��d���]���>��?h5��A����J����Q_�нD�*��.���^�H�B����W�ߩ[�M����\8y�l��uT�5��6�H�I،���0M�ci�7|�x\u�YO�N,&mR�0��m��U~��
��E�)S��zU'�����E.><�y����>���x.��w0X\�f��:`\lY㇩o�흓��h��O�	�բ�7��G�����qc�E���@aܯ1��!ݼ��������ezh��-#J~��l��mRKL*>��Z�ڦ�4c6�%�<�8s�H��*
%j9�''��*��(�Wsbb�X9|P�i�ҚX��wb+N�z|2��ʕj�ڤI:v2��73�0]����q�s!�Wz�yU�8�K"�S��uVz���|�c�E�R�
j�4y\|�cG�[յ���P�����BGR�p��� 3fp�d�t&u��,�;c�@[J\��,<q��ۍx��]�|�]�{�λM�����
 r+7fR=���
��I��������v�'�}�p��=����)�I��}�S�����&�D-UM�ӪvڲZdR��Ω��H׻��u�A����'�"����̑��t+��e����P�lΩw@����v/�.�����ֿq	JV})�
�4�r�
ް���LR.Y/T���M�-I[{�e̺W�my뭞1��)_�*�>����a�����\��4ڲ��G�llq�|R>���<��O ��M��d%-`���k�o���ިD�/��������E��p��s� $S��T{���+��!e��,�콡��oD�|������Gl���+v�}�y���)yw|�y�W���r
�zK6��;P��7�j��3�(zhD�E���r,���y���qc�i�*&f�!�C�r�p���.�?k�U��;کQ �����pp� �xo�;�=ض0�]�w����9�� @���;Ӎ��7�M�T���Y�n��r#{���˥���N�<���:利��Mۑ�̱�P���e��oR<#�տ���;ڶn�䯷�S�r�h=G��7�L�k҅��ި!3���	T�c%O%.U<MXIO�h�7&d��x��h����6�*es�%&q`��H�<:���!�f3A;ejF�^՟�<����a��Qg%��T�kUȬ.d�mS���d��l .ž��!�+ĵ@�B��҇$����o޳�2��J���0DF��R=�a^z��a���v��.#��������6���q�{FK}�����aLiNM�p���Y���n���+�gAA�����B�ܞվC�ո�m���p�⺫�G3���2��?g�<V�ғR���[��!;��xE��q�T�Kt�ם���7ji˪����3�Ucm�����B_��:g\=�S�������)�z8�i�I�;O�v:��˂lc�צ~"%`X1Z[���>j�[�a�X���]��|c�{�ޯy�iO��������0U����n����Ķ�	��v��Z�s�_���jx�]l?��KB�m^q�7u�p��Q��L�VZ'HW��}�0� >ݿƉP�����r�l��2�2`��O��g[6,�������i�Z�~�s��-�ga�\���x0y�Cts��/	�/1�]o��)x�ϝ'?i��` �������mn�	M>=_�3e�v����)���jۧU[H�����������6��w�U��-^&V��B��Q�m���q��S�7�x��^��;��Zx{�� �h�y\���čGR�.�%U��X^<��k�^��wX��t�M��ȳ�t�a讅��<���b7\׈�]�r�t-wo*���J�nV�Ǧ����%�V"*�Us⧣iX:rF��1T��ָ����rZq�Wg�Б  ��2{���7)��:��hat��zݣf�d���{�~:�8CJ6��1�>�=�����-� :	���g���AB�q��K�Ҵ0`�8[�W��IDJ��d=��a������	��\��r�D���J.���v���i�������3ri����g$C�R]>��ε�K?L��_B��,���.�#�aa�6U[Q"Zڣ�B����@⵵���sL1"��v�U������
u�L�������~0~OJj�e3'�j#\���7��!�'C�u��t�H���{?��τ�-�_2a��H�|��j���t����+SAm���g�������L��B�?��
�]'���HsK������z�۸ꆆt���{�C�C΃���ĄUYY)�qI:=���Ͳ���/�)�O2��
�_��+���?�
/��������쬠������+�z$�R\J������~�f�J&N�&��?��L����ה������<񎋋{����ϟ?�K�Q������o��_��צMFJ��Ƿ��54�588���������������I���ӭ���Y����< D�P_600P@Mmr�hݵT���W1Zfcaَ�Zw��۳}_fI�T�����t���W
�	��%%젢�gdЉ��A/���q��_d������d�s��`//���Fa/8xy_b��+!�韮�����CU�1M��6��~Pp����V,��蘒���ؙ�h�qy>GI.�oMk5�H����*�������tu��u%�u���3ps�|�z������y���̧��J�iii=�)��%��]�U�m1}����11$,,,o��dee������ζ�x;�'&T�ܽ+hbb���n��۴+����67���h����8�2�����BBB��RR�_�^�AG����#�����QZ/'��䥥��������5���NKK�i4g���srr����G�к,�UޠaOO����20b�Ѐ,���Ǡ)�Hll,����l�	��EES�kkt\�ƣe���߆��RRR���yx�PQQ��FJ�v!�Z[��)ıa���v��RC��㨵�,�Y¬�#@kA---Mư�'�����yxx�vV���K���=Ʉ�cXJZ��ׯ_�����{�!/���!;v��=���S��i�t�I�lXX =��Z�ÝU��	ٙY��4}�.����ڭ���k�<���1|1�;�?RR�{���\Y���n+���65�:<<\}u���	Z��Ey�O@�v������2k�N'L�90���ۻ�ׯ{ E�������_}}��������A���(�2���u_�nD�VP-�Uxll�#���BV�?*ŕh�v1��@�pNo H��Ϸ�l}oӎ��e��T���HK�#p�]3a��#yX9���W��QIe��\]]s��J�42��ۣ��e�@��:�@����^�@=���>h����N��U��!!�
ڐ��!��!�l���E�,����o���	�?�3����T�56����{HB�����n��iim_Y1���OD��{�g�HYEZ_Ldfa���Y.�/++��ۘ6;@�Q���+�3V�oml�C!~ [r�B����|H��A��H�.��2������ /C!��5,,,0�"�󑭥��@� �)-�FK�ή����:�u�+,d����}������������Tj�d��JK9��G����n߆F��j	.��P'�s�v>X|HD$a��Y%0;?�8�^�OL�XZ^&h"�q,��^�t�y�r��kbb�|qv+
�Ȗ��l���`���>��� <6�qŕ�s��ǿ\��gDD �PAA���E>���x���E��$vƪ�틽 '��ň����q����!111��<
`��h@8 �)q��w�����yX%(�����S9`>DT֫C8DDDf3�~��%�\�_��ZY�h���x���V1].�#��nկ���l��������5Q���7"�4շ�zE:�n5ut�������B*W��N����--��L��6Pd����L��FA�$ �
�.�Ä\�t�����֬�zto�ژSF��Y��cqY�|�M�� ���nܸ1o��=3����A�PL���c\�3x��|G�or�3g��\Xht4���WM�u�!��~��^A8�l��
�t��ƈEǭѿ\b��Sd4���z �08���r���Bө���˘t�4��y󦠨��:|�nZY���-&�Z�@gg=���Elq G�4
�Aap)(��:R+�d>�<���Xe[i���&�Tl�}gu�=�� 1�nSMT1^����Q�����ά���~�Fo�Ӊ���X-�yT�[�����Mf9�uk�T�ah�AA!I(W
t��\�~����2�ؖ�!0�Fo�,�W%�+��lE&��B>��;;֙$�_j��Z4s���JN���/r�&M���Q2�d98<��"vK���5]�8%���h�����b�ń  )�UN:�";�����"R��$�����B�Ķ�l��o��l�5�v�OH]S�|Q�o�xB�ݸd�kJz��=ZEpc�j�0�����?���g����@$vhHRR�s�~dB��挗�倨^?���p���\��j;��i	{�Hv3Rt"Nl0��6*oX#�W������f��xnf	� �")��Ҕ;U�����%.e�F�x�J��,�rR(��C �@����{P�82B����$�AzȐ?|�TT�P�E��G <�!#$d7��s�9��.g��4��c�� X�sA���6�92B�˽)��
�"��|��?AWf��}�J3�1;�cd�ƀ�oCO�ۮ����K^W�
�/�W�@b7����#V�ǉ�$#�}��l�+@����S+P"8�l|�\	� 33�⇻�YYY�Q�=�bttcQ����7zT�i�v��κo���ϔ�$Ν1ӗ]L����l�<���jH�m��s���Ў$IDLA�|SSS	�����@ ��J.b�t>Z���'����@�b>�q��l!�.D�i����]�S�B$���D������*do��������{�g���K�߉m졋E" ��^�����.�a��}�X!-PMVN��H� Y(x�?��x�q�-�l�0qJw��%٦�rA\�_�Ft.<7�o�䪀J*Z����nj�@�ؔzG4hB�Q��@��ç}���x�߶��C��+�V� ��I�����x�?%�}J�۹.�'��^6�' *�*�e)���h	/@<W:��A���I��K�Ni
�r�B�d�Z����f����B��t��E+q�����%�u��*ޱ��������zw,�3Wn�ȇB�-&E�ƵH�]�y���bD��:�GXX�%4� ��W��@�DbC ��0�=�N�~/  @DJ��?#�����{O�qŏ���D=}}pT�{��H]2@k/��'�#�A[�5P������7��A`6o��O̿��?i:���RYB��oee5b7A29��c%�@H��\ۨ�;���.�
ظ�Ȧ �qK�����Gj\�Z���!Q�c�q��|G����eJO��>%�������r�U�Oۉ�7�@�%"5��^넧�<�Ӕ�?p����Y�BSj3q�/!z��,��722 f�>�8�5`w�]�=^>�9+oee"ƐI9j/�d�q�4�f}�*تjץ�,���"�DW�|R��J��������7��{g��7�R;4�UQ�O�+ǋI�
Λk��Jh��f���%�\�Դ�I��O����Q("�'�Rח�%!�S}����\��{҉�W�.W�~;*1�ˉ�b�s%��d=*>>�ǔa|.U�h_�?:�755���5Ά����>2�?vV,�zo7tT~�}�엪!��V�1O��~^���.�Ls0O+�|VԌP��&usz� 5-m �."�����u q�$@���A����4L. p߽�dɞc�{��#�:!�	ӌ1������OT=��?$��`�?"ff��}z�u��Ua�e�PJޫ��f�+/Z �F�Y�
� �zB*����X�u��펂*<�����$�������ԏ�bN���;b�5<����g�RXs�~�-!e��(����'''��2�UX��&6�AL'g"4r����>c� �kl,�:���4��A���^E[KG�c��X����P���R��~����K�+8v2���kn!i��Y���2�?n3�q�{q�{q�g��{�IQ���d;���8�*_��`���TV�iR�P��(r�Yx�"��7�Hʨ$��Ր�����:*a�y�{wFx�������v���^y��f����< �H����7�*출��Q������ޘ>_�t) �Hӵ��NN��й�t����0������H/_�g��&rvP'&�;Y�`��&l����Xd��8�����`�` ������d�+IIY��&`�SҨ�n�&���r��IS���k�V�1KG��hV�l�+�9��M���,t�q�����:��8���Ef��������ꪓ���D"�30���GԛSCF������!:\���'��9}Osb�\�����@�ܗ9��_�sO�{1@6��$�p.���=?%�Ӻ�[�RR���+a�0v�5\?��ݟ.Χǻ���]��־����A6��@�Q	Z��FЖP}������Jx�<ռ��\P�������c�m���`�.��������+ww�m�ݶ�v�[0R�M7�=�|����11.�pZ��4��q�&<���p&H^��������l�C���1D�8������o����AÁ����j������QRR�MR5���9d2h'~{OKJ����ȷ��۷�Н V�Ag�FC�6f��l�_(�d���u�=w�0��d��h��f��o�'��߂m�b8��v%��bc;�?�������l��縒�o\���xy�_��ۃ�t��������&g�//.�1��<L������;-\�2h�~C�P!o��in_�=L^R�д�t
���k��C��P-��S��Kq5Ȑ�	WTVg��d~�ǠR�d�����؆|q:;��:є���}�`�5�)��k��#~4�>}����퍍���l�QX��p�I�ËA
ak]��ޯw	�nvo��ת�Df�E}ct�l���9R�sZ��XvKl�2u����Mp��I��xZ2�jWP6(�m1�n��t�rw����h/i��7�)�������o�6yBOS7�+�,������TT�!�˪��!L�U�lnm�T��T�d��������׊�HI%H�,���<��( p�;nǯ���8�J�=9�^�=�'=*`�a����Vb�Je��ὸ�#>�A!�܁qh؀-1 �����f,H��h<=<N�DNTA����HquRJ����;��v㛱Ľ��w8�Z�eV�!!ɀ��n�� bCU7i���q����hI��Օ~�W��=t OQ�W�	�V�����cqQ�3��~ Yє&��e8υ� ���:zqee$,(h���������xu�������&�.Q�_�vy�� gV��t՝�0�����ifE�0@�_�����;�L�W��<?i�>�Lp�bu$I�ˢ�9����;��o����́(t�B��`jT@�Ò�0��ls��ՁSY��"� �f�u:�V�
�W��w�|	�������C�t������恶�Ʒ}	WWW�6�-L��
�S�Ӈ v�m|�_�,^s�$�X���xy�!,������PP�4��hֵIsS�oHʣ�|�Y���-(¸L*�z��M�Rʆcvy���p�䒯�r �����Nz�{�n�D'�f�6Yi��i��R��[dÙ-��gp��>�/\���1��;��c�1\��y,jb�>l�F�y��nk��5i�g�v��j��f�u����N�P��Y~��U�Г��N�<̉ezg����Ymllܬ�F�K�1����Pu�Y�u�ǂ��y]�r���&(�������_� ͏����O��I7K�<���G��N��H	�$,8R4���h�ٴw%}|�y��3��b������q��[I�2��P��4Y*!D��k�2kc�ne�HDbH��%c+ً��3�g�>_���3���׽1�<�sy<�s^�3�w~D�4��h�ĭz}M�x�2�����4�8f���w���8��3a���m�H�F��t�_����xtz(JK�͍H�P��e�ίc�`�?�w �,��'�̘T�\I+�Ǳ�w�Z�N���>��m�R�`^�4k�hR�Vi�R4��"�4�6�[�B�RHܞDD�=�kRXmS�Y�������8����d5�/�u�%�Ƕ}7�_�\�$��>�ӽ8�|e4�\S#j�R�A��)�� ��6]s1Zk�֪��^y����&&eQ�\<O�H{��F�R_ig��Nt���Q�w�H�-@^*��OZjϐG13U��˔���4"_"����τ�M�G�s9�J��R���:s���M�D��r����=87��\���g��������pj���r8]�5�=��=�3g���IV*�F筥T�\m�SD ̮A�����T<���\�[�=�*
~���1�V}��D%Y��g�
獩(��lCb��H�~��2S�H��Щ�����]�����)
Y�Vtз��e~���B�$� +�7��w�r�[�|���?�̷�	�.��F�2� �3+Ay&&&��q�*W�F"�uv��ފ�e�D_H�,IE��^�����\���'�\��k�O���N}`omkK�Gz���a���9�X��ˆes�ː];k�{Y�0�w�'�ϸ�~��*�L�nQSW�^u�lŀ�;�+�����%���>�8����y�E<���O���=�Z�m��NM�T0jeśM��4�*���a����H���x'�>��f��BU��B�1��4W�����o/oc��g��
]F�Y��4^�J�o�l�������g'7z�TKSp����O�\cD�mj+}�'����)c��q�J;���CƆ�0h�c��!����L$R�.R@�|}i<7�_^�C�N�M�H���n{WL/��@�d���s��f[��FN�CG6عkW���kFJ�K�l.`���_}f���~�W���ȼ��0��uH�/�qp�$SO׷��)�}(�w���z�
?�}��#M�fb��<�g��`�2jaϚ�}2DY�d��1I����s�o�&�K=�T�7&���`]�<��S����� �.��@�z(���U�<4���F�71C��鈴O��� i�?�������o�6��'���<��s a�6�k���A�e��D9C��{6�T�c�#���Z#:�`�onv��SO
������L�|	�y���(^a��v����1��������(
U��
���*QΫ�5�Y�Dk��F1���<����;���5<;�F�7k�R�eJ~��* vuuU���=��i��i�������UK��J1v2���cTMM����ЇE#�)��*���%�� �ԩ/�L�˛
P	��t����6a���p;7O��533�rqz���~�f��k2�|#�J����ޞ������5�pQ0�"��{�9�G>N��l@��1��V��??�J�;�Nմ��">��׶�$�;�{6�o���kvo��G	E}k7 �@ΰn��hr:�.y����vi�P99��Q���-rqȞ�8���|�����o̽B ����:�rKF�����>�&��s�A�7�.!n|��N�Q\g3+]� )A���� lP3k� Y��$��Ԣ�.ʂօ��lq|(�`�4ȸ�J��p��:ُ!۩�Nmmm�>��_�e�n��P�~l���g#(Q�O�>�k
��eo!T��*��z���(��G/^�S��\��i�q�*��<e�R56�d\�o}E�6QSS�kM#sn��|��5�t�$V3I��<�%�Gzz�
���w��V&������ˁ���G���I����F���Ȝ�c�N}D�>�  Ѥ0�P�!+j��5ccљ�殦�Ǚh�6��b)����0'��'�so�
����/�]Ϟ=+����և�!��%j���F1�e�;��!Z8߲��6E�C1�m��C� �����̑��h�r�#_\��xV]�*��jm���E�j���S���u��Y�H�W�5�秉������X]0a�P����8<4T\��7u�f*۶��Q�l��՚�A�"G=����Y�������(�I����OB2�q|�k�7m��45�=#Z����ː�x ��vv;K���_% j\�P'=��tܸ�:=*�<^�dّyc쌼}a�X��טV�-�l;�rY��]����s�t��'�O��ݼ�m�j�d�왟�fU��A+v˵ �h���O���b�a?~��I[����.�x��D��⳶�������ަz�.4|��0�B�|���v
��0,���X#����&���f���p�ib1��B=`V�P�_-)*�?�>�+��2������a�w8��	�g}hf��۫��m��O�2I���sJ�����QBZ�M?��h/���rJ~�E[�κ�4��������'�m>�^v}�kԛ^^u��隚:�yz�H�IeK,����ok�Q��`Ȣ���Z9��_���>�H� :�M-�B�WV������W�DЮ�8�Kt�X��G��/��5�>h�Ħ��$�oBK���(���N�|������BX���DWwa��tB{�e�CC����Os�^�O�� ($��'�!��o��O�U�����{Ё`蟷�%(e�����r�6���S��{��%�3#����5a��ZJ���v�!f���1T�PU�U�u]�Əq��F�(1���x���.^vm�qvaA( 8�7��OMW2�酟��0���3�9VWW�ἜsW�z��{�Jۻ�����Y� fEc�c��j�ܫ",$��-\��FK�tuq( \
t���A�%s��/<�rT�<�����z@�j���V�lcmpo�O�>>�7�|�|Ｌ���v��ɽO�r�榦k|�����:9�uwq�y�}����/PTB}���^ qOV`ۖ� ���	�����퍌G&3Fo{z T��X_����漕U��s�a2gNu��>��l:�P������<h�uC�Omv��m�ܜ�X���ma���1��y��/jX���R0_qL�(�t
�!��ý��au���X�1.�:s����vq�����h#n�˔��bc8Z~T�j�+�x��-���y�`�	% <�I|�O=G�1���	���2�#5�t�f�m�3��W�@IG�d�+��~�W��"�<�Z�e/K��S�|��. ����*,.��D����K�姌��)MrB̇��d�q`��ƴ<;e��㳓��;�*S/EY���2gJ'T���,,gȢ���S� ]H������#��{6M��1:6VHaKjW��;(m��JQ�����7�� ��@���被n�ɳD�&�H~^����u�p��e-["����|P�S��Ah��t��Y�q�B��
\��Ŭ>���,w�������<]?�/	���8fD�Ѿ|�!�k�����w���O����O~�����hoWur�O�$�o5'������#˫KKK��C��>*J�G����<E��h���@W��/��h#��^:�<�9y��{?��^ڸ��R	B�s(��L8�e����x��~q����\74\���6��b����yR��"19��ܵ-�N0Ѫ;n�z�m���*Y�.2��������S���|1��%�����	";�y���y[�J_����{�,N �~�.���3?&�����ud�x��s4ٰ � nkg�D��o4�ܠ�xf�4�W �]�i�o �t�Y��`(��`o]�ZT4�vW�^;�$��:tC%��V��EE��([ܯB6�#̔+D��,*����j#_�f*�^����_cS��S�;"��[�@%��_��ŸFU��6���3�$$`������H�v�f��5pc�����g��
E�h+O<����Pm�4�H�7F[�`ᴐ' g����Ϧ��+J��İ�R��T�:��~ƅC�`z�U���9��|� �C���g?�"˵u�z]ʁ��H@��)a3k�� 9y��g	�\��uc���H��W-䷉��'h���y1�DU,��a�?��m?5<23'g~V���]gOլ\����Q,y����|��V��Ͽb<����Ν;� n�.r��Ç{l���ss.��	)��;�O%݂�=nR�N+7��%�����@Z��$���Lz%�򎓝k���c��S�~d��&�PX���]��fy��#��h��;�����O2<�+rL��j�=����kܶG9ܵ�Ԍ4,�O��Rn4#*�~�^���
���D�ieS�����܅`�n��5���Yߛ�7�7Ҕ��;��^�����_�d��O�<R�?�R	�P�}c�&ƅP=H:�A:P4R��v���т��J�1&��]�%M��jb"��E�K#\��c<>/�v	C����k&���BC��?-�,g���rbGm���c�w���v\\���=��v�<#C$��-��U��y<�;��ˊ�����m�>77��qc��߷s5*x���
aF��,Ot�X�:1�x�:R刬��
ޭ����_dѪ����q�e����׎#�ra��eD��U1���qy�l*E����Xk��L�ɫ׮���[�x<��Q��l��֯UA�I6�ϛ��ǘ���w��#���,��㾇�i���
"�������%�"�Ǹc'l��JI��2��n��q�BU�V�Y%�E�7]d޸ߙ�����Y�N�b�	�/_��d:PDH��u���e�����@���w~���� ^�G�l���E���ۜcn�P ߄~h��2�
g���NX��H�%���M��rU��s,-�T&�"�C&�?�lQ�lN������_���m�!EX��Y��rb��rK�E��k�V�����=J��)n��e�1Kii��89�B\͛��&�������o�v!��sc�J�5���M�\�ĭ�ׇ�^5,<������DWi���S5\�X��w���.�}I͆��111nn_�2`�~�}O�MI-<!+3�1��鴐� �O�2j��%-�f]� �ʩ�f��D�Dʛ7W�/�m����
�V���|�*��`��<k��ړ�и	sp�xG�-�x�%�5�V���WG#��J�����0
��K>��7��i�ܘ{/"����ҁã-){&�ʖ3`_bCC�:1%%E�dq�3Xݖ�y���P�׌���F���m�����k��'����=<�7��a|E^SJ��3�I���2����~�WKu��ڬ��wbI�B��vz��+���`%�`~����d�]��8ت.ޡ���TpL�uI�v�5,Z3<T5���{`P�!s��JS��o2E�{f����?�������K�z��4����k�N�e��",�%��~��2�`��7���V$1*�A�������_��Nbb���ai�{d,ha��p�G� �q���kVa�3��%�a�Ex�P��|MQ�������S:P o�I7,/�+i��&K�Ƒ5�f���_�� �m&md�Y��W�N �J��X�N��l�v�����@�,p�$�VVV׮]{A��ຉ�Փk��*�����[+"ҭ� (�
��ajf����r��ګ�إ@�ځ��T*������d?r� ��Nt�[U��"����C>C\��L��Y_=�ptQݗ�eЪ�[�
���:��l��[��<I�-4������,�:�;a�W�x���x';2A:d���09�	PT!k����T]��&��$� �?�<:���7�8�ک���6?��2�#���ES�/����5�k#e��];w�� ӑS�h����Wd�����<��u��:�yt+??����j�����t6b�5�� %�$0���x!�a�O"~��k^Q��j�%ٺ1�������)� .��Ǐ���g����:��r�F�s��d ��E&%m<��iql��V���/Rn�ğ)�B��FZ�*�����'y�N�U����Pc'K�spT��.ZƂٷ>=K�K�Ka䡫
=��I����CV~�4�
:��E=꛵C�#�f���'s��Q��P���ty;�%�ԛ�6����� Rlͳ���un���P�یx<~vUO�hZZ}뫓����)�e��8��M7�}�|�E�S[�����	42�� ��򭦄W���6'�RZF��̓)0�9ҡ&gP�6��?;��I�=ʥ@�Ʌ�S������%e7 �1m�c�V2�����G2�� ���̝���2IH
����̈�T$���,|$��G�y��='����C�$�yT-+�8dE�UF�܄Q5A�ֶ��X�Z���	o��wfW���sP��g8n�CI�,�DyV�i;V����k7n��%�H���EB6�Y��̙�kE���������� 1z�/����Xc0�<[̼�����dJ���	���q�^��jb�hJ�[֧21:���ڃ[1��jVonc����M$��A#���$Q���mp����W�n F����n����=`�e7�|g�:ۂ�������y���x��Űz���s� 	5(�d��y.8q� Td�%�8�t���}�T��W��UTT ��eff6�ã��W���HÅ (G{z��� �}�i�L��ɕ+/^�H��v��~���	^�m� �Mo����[�����<��2
�kG�s�G��iy�� #Ҟ\��T|�F�2@���S�13�Z�VZj�l9�����ya��|+��0^�n�I�y_&Y]\\��я1���~=�G�b�(]]^pC�F����l���?�!�4UC$o�xjPZ������N�w��r 	����d�djNN���v� ����:w�X��ٟ����T���G��3�L�{��J�H��uXm��G���V&m�O����B�9zR��,���?�]������(#��]r��n�-�V�}��:�!~���fr:�,���`>��4����8)i2�Bu󘕆�o��Y��Gɻ\9-x;���#Qj�0V���ham{`{Gǝ���)(�OOOZ'D�C~'�]߷�٦Rq��O��e�p��0[Ȥ`T�K\���9�� /�p�j�W))����K8*y�V�(�t��5���5�����/o%����6l�[ ���ȏ�Թ�2H�_w�;�LM�G��.X[�T��0W�j��u�*�h��+�XYQtW��Uj`2����E����@��[�M��j��i����?R=w.�?�x�˩)�f����Ic�k�.��s8*LRy�$�m�ޫ�H�~��8#��߱���ׯ�+�����ǭ�q��5�������,�<�S��5#3�d��̞���!�޹S�N��'~�t3���Y��2�����uq��J�,#�s׶4���]:q�D�ZW�J���toy3Ԝ��ߠ���1�PZ͈EI��0"r��-?���L7�_<�������J��/�vP�d!@�q�D��"D��9���<g�����U��]�1Ӣ�?��5㮍|����zO ��A[��,tW��i~��?
��8F�{�}���ȸdm�t�I���
]2K���g�x���R�S�+[�к�d$���r`�0����{�E1�I{x=��b�E˫�]�.rJ�W��rB�hok{{�d~�d��(
�9:�^*2�<$znv��u�C�szQ���K��	(m��ã�h�� ��.n�S��_�t��khx����u�P��" �ko�B3i�O"�˼٣�2��R�H�Ѵɻ��`��v���|YZ\]*���<�ӷm�[~���0�vf��V�"���֠6��Q~%:�*)q�z� y��]��u��̼L�pe��z�X7'� /��E����#.G絠�P��'D����0I\S �4<?B�J�TRP�K�������F(��5^�tY�����|�m��/�_O�P�TR�0�ͼ/�������cq�HkE�Z���z/���T(�5��'�4�]���޿q���Ƿ0u�!ވu%��V�ʬ����"�D�S���q�K�J��]a���]~8ܼ��(22���w۶n�oj�lR�'����9�=��އ�y|Pt?mN,%A���V3nm6�ҧ���� [���O�Z'�2���j�r2.��lkk�joo�'p�G�E@W�6?"�y��Z�F%~�7 :��!�����ф��I"US�h��0�t�wX��T$It�	��s�Nt�dbb
�ˢ�L珁����8B��@�Ώ��H���EFFƊv,� ���Js�ː/Z5c��Y�
j32���.%*���#���_/E|�"
����*��33�3�nRG�|8N����V��Ĩ(�ߡ�ӛ�u����׊E��w5A���K�VI�{�:�|F��������rH��Y��D�L&$�C�rJ���;��X<^������� �_�5.�z��S<���Uh���y����ge�N_�.�}���d����JC f��8�VV����*�z�E��Z�f��[�?'dG����WRS�dr�?kֳe�H�э�t�B� ��C�E@�Vg
���l��^�"[D��-�#��#�7��
"+YOWIiIA\.��l�6�n^R�G ��"�{���S��Cm��a�ho$����Uc�=��j���d^'o'�'!J������Ĉw܅�r7�9A�D��Ob��7�S��b�r�`�!����߄�����*u�B�-X��<����[3��_�p$A�-���%���T����߿�wm�N4R�P��̽%�T:u�X!�Z(���4�}D|�0�����[��I�3���n���g����؜ȁ<"��&���������v��0�k�{�؛kt+���L�O%�-6 �n��v��MD�$��+�=2��\n�<�XeS(�(Z\\�Gy����)�$pӤڑ���/lI��&tD�"����7����tGv�/��!��-'��?��ӕr�.񗾾~o��0=&c��>ܔ�:l�8�N�8Jb��L��H���;;�3wU�t�p���,��L�q�c2��b�*'3�Tme�?��o�F*�����~b��|t���׬�	]��~����\]�}�zK�W�Nxj�ߣ�O#����e���������t�>�*�:���pi���į�`�j��w+�>�l�y���=_�-s�n	{��N�'���p�������=(�rIA�
��wT�v��K�<ʀu��P�e��ߌ�0�����Ţ���nAgG3+�!�R>���A��g�!J��Dhz|�����S7d�|��,�)+{.���G�*�+���u��9���L�g�X-�"H30�(}at��K|d�����9�M��{˥�:k�/8��2s�T|l�?��V����]��������8+]- P�4��*bӕ�5P���Twz�]S��X����a�s���"��G�����|H�2]�b<j��$sJ�u����
rV������_�
�i��������Gި���׸ty+���7f��C�ִ d�ݩTѽ�#5�S{��o���IX?��ԖJ
5�'L���O#�,�Mܿn�S1i;�ѭ]f�!Wݖ�>����7,�gr/��y���T4{����"��B7����D�rI�#i)V^Ia����Leӽ ��թb�	!|F�1IB>)b#ǚG�6_����g;~�|B��4y7�E�~L6��R�󱉒���Ns��ň
w��c���}��N���8��Na���b����.�_\	R�O�KDߦ��,p��Ɵ�lM@�Ո*0��EDD��H�6��6����8r��zP:""�|am��V�`�׎C�{��8�f��jok�{�����W뎃�{5)���!ؕ��Ʉ��b+r2F:���R�Vzt�ܼh���R�9�{e�dEy�`�ϭ�m���t�Z�����p��a�ӧ(ss�,@l��Lw9%%;}4k�+�9�Wi8� ���XsT5y75o	#�y�Y����}F��r<y�$"�冇�����_�b�M?0����-�k%����6Z�v��c�_&�	%��P�Ge?H�68(��ݱ�9���R�l���ދ%����⛶�M�.����]n�o0d����+���S]S��V�P۰��\�Z��8���vF:0�7Bm�Z�d9�U�VY��c6�\|܇Q�a��T�O����^�L�,��.F��S��z�q
vA�����].�,^iwo�ڥ毎?/�Q$��7�R�G���9��y���P�8�����[1��^I���۸�3��LKRR�w��f��fs���x���5�~��OcgD��3�r����۷�.xe��ҽ����hr���۷�>�����-��d�{��P�ڑi���x�b��9:b�i>׸o�ԕ�/}���h�v�{�e��wiS�Έ�w��e>;s�y }��@V�C�ܮq��M�B$�����9��K㓲�'��Z5mt7�Ȱ�D��p�]�'�{��e�v���A�Сsm�;hf� 5�(X"N��U^ /����C�ꃈ� :o��=rFH��w�5��^챍��$H�$���L��u��������'1� ��A�����
�l�l7�%�~i򓄄���e�e&�����O\��i����pllR���r������亽܈�N���}m��4:z���;vިʋߒ�_etc�#
I��$!Gl6�3/ڇ�M'�|\?z$���h��[�������9R���e5+�k�`i���!���_Z���4��S��8i&�ӟ ($D
�Ç�y�EOE5���ngMh�1�0��*�H�+��40�',A���k��7/K/�CF�իW7QʊH�~�����,��4k}��ݻ�NMCc������e{D��9R� n��c̛�N�#G��]�V��/(,,����s�M,����i�X4�lиGg����B���!UA�5v���Bcjj�:t�/w��y�(�Y_;d)�|c��޽����AHH���yO+�&��ą�KBZ�х�� ����b�Y}Nl#������8A�O��!��v+�V��zU?]���]���q�QQQ�PZ.+�����;�<�}Sa$)-ݶ���- *��+��02giɓzO,�(�<�����c5d�����Tf�SoU�>��^;�JII}��L_ ������kjv��:L�Y���z�{{�SC�=oĈy7Դ(]�4��)�`��ꊐ=�+K�0f�~+�bW�߾HF���GP���5��q`�)ZC�dΝ��ՠ��U�aE����E
D���> �����i~P�a�^9n7E��qT�2F�����%�G�86�V@lKj�A�:���w;V�����Q���j&�NƷf�ut����v� ����Q�ƌ�o}Dqpp��C��MǸ��@�9!#��&@gWWR(�r.>���fkM��b�y� ]"ȿ�P��?��oɉ��n��5���I.Q��y�e���7��
E�8&f~?2n4/�=F�5.,�]�8Ti�4�kj��������H��߻wo
�"��x������������ʪ���b�̢w����qjx���w��.NT�~N���tD��+1�����c���I)*����S��xl|��c�;͠��duy�;��kUP{���i*��-��W��~H &�\��H����'N�Rsqy��� �7��Z����B��4���^�t���F��0�[����ȏ��r��t |�'m������[O�"E���E*����(!-��\�n��+r�Y�!�|�.�SVV������w���m�,j	�g�qp�hA� �*��t����ƫB�`�Ksss� K�.`0������`c�/+ڑ#�V�����)	p�����'�j\d��X�KKϲF�"a|�t���Φ�G<&�
ZJ{z��I�N&�OCC�3�!{�����$��t���\$ާ+(�/��cs����g�!	$a�Q���22n	=�NM�X�g�؋��E`�
��כq��������PkcE!��<����b}t���!,A���k�ܹ3�'����	�S,�����'���<9��b��ǧN�jjj	8����a'�Y���{��in��E] ��-�L��:���#�-��"}��m��OZ}�W��VQjLJ����ϥ;����e�r�Kum�:p]HS�\�VE,���h��(��vgΛ�w t(������k���Y@
����H��!Kx-�:4G{$P+��3�,��ߟ� E�n+�H̯
ڣ�i�0a���DD*�����DB�"��~�����@&j��}���Qd��o޼y2,�Ғ,����/e�ŕJ�};����
�!)����dv4l�Q��>x��_a
����$eV�/��\��b���jԃ�Й��Z��tj�}
|�����zIU�Ȑ�E�?^�J�<8�OFVE��
0��{�וR�������y��%�7��{���e���K��%O�%F(�?9y�ٗ)Co+�WUޕ��&�tkC���/�jb�'. 0��@8A�f9)#���S�S�("0.�k�HKN>���M���n!((�+��߂���횶vF�5�8���Y ��{Q����4w�ǚx^J�]�����?�ܤ���o.�L�����2�`)$ pB����y)i������������N��r4��x5X
Z�٣ȫ(�T)��em..��c��6�>���O;>�u-�SّR��p�o���!ix;����ֶ�~ z�I(I�O,�!>�����WcD�@q���O��"ty�����g�n������U�[�˗�1b��g��Y��Б��Mr�֊{�1/^�O�p!��؊U\_����yd��c�������3�?�"�L)�s�������ove�[˂���g���R��s����GFG�>2G�9y��,��8�u6vv���aV�������fl��o�`	������_D�N������USq��C�bb1#�^����
.�z��`mc��|}-��4
&4>��$���̢Xĝ�<�� ��8�&�}hp�W{����U[;;;��V��B�Z�K����\�.S	m؀�"m���Oq5?�uZ��u��^ּ��4�k�F��*>�VA��GC\rqqዾ�<yO+d�r?�_�JQ��1t(�s\���*�,�W*�gϞ\~�(3��,s{��LW����9I\Lw�7nF�o)�t���_�PL�E�m**ߚ�|!���̋#����3��Yh 3�|�0 Flg�5�7�wre���DZN�f�n�t�B@I�̾�%~���5�;:�~{J�;w�w��λL�;O~,ZM����c�:{h�X��ė��� ���sʆ4��	@�R����8�<	��C�U-,RVF��2��JY�\%�.:;�_��iЭX�qICc_���M=.��g��`=|��CjzzÃ�"ŧ�{Q��}�'}���Z�����������	]ho7����o�m���hvm}m5!g�j��ٸ�z_n�q��/�!L���l�;uq�y����G8�\&�Ŷ���R��U��N�ɜ��x�?u�\9��X�5�n�Ժ�sQ���Z�L���U���ڭ�"��O�KN�,j��9������?��.I�z������6<�����9Y�`R�����O���64I���vmxc^VXX8	zh��L�Wg�H-�j2�-����!5�%���G�0�������d� 4���5�k���5��~o6��퐼�{�\�a�4C���NL�Q�5`cM�gy#>��h%���B�U�a憎�ܥ��;��3u���B�r.,�`��/vNc��*:���[�1����g�e�:�B�-��W#��La�l�փ�е��*e�K��X(�YD1�Y߻x}w��6�'Q4�p c�H��/�w�o��f�?��c��)��W��Xm<ӧx��4��]���mjI�B
���ĴN1���w�@C��4r�znPZZz8��w��ho$�Ы���P�b��C�/W�~+ME����毎����j�\�����t/��Ǚ�N��}e��C�_���LJNV�I��~�,��� �������u;j�<�t|ˡ��8�-��. ����i�_��y�jj>&9ď�2T�!8,|��Dk3r�̋/�vl�N��hD�9��x�ۻ�����OmB��e�r�tu�6�E�u?���xP ���wy$�.׹eWhj���>dNs�;�c����Nq���W�z��� o�>�����]����4X�֣`J��]���T��ϖ�֝����œ����.�_��̀3��u���h^�MJW�9�������_�.�� pw��𓗑w��WI�-746�&y7�O��9�O�C'ΫU��8�����fh|��6C�4�i���8N2�j�K��J����u+�{�߲�H�guh��ДC~�����ŚC.���qMO�
hU�_ޘ�)�]�3^���'��:cù�L ��&�h�c��+ĕ�F�pJ]E\Ԓk��S*RՒ��V^n�,E�4�K�����Y|�	fY�`��+W��o�" 
���JYfa���!���G�(<?��u�~[l�N9ԟ�n�xy����!j��&�"��MO?�]�W1C��[�$���>K�f/�����AJy[hߓ�w4	�!�K�h^Gq�� #��O5�����c	�:�G��s�[����xYzv�'"��7-,���\�`�H{��� t�����e�};m��ݸ��{Q���"���v��w{�RՀ��@��gfBzz�E;�h�*^��7�}e��4��#<^y��4d����V�Ϥ��X.� �������k�3J��Ϥl}nȝ|e�E�Y|nY|�0ڍ���'��{������������N��f�.#Me�@J��-�͑��W�k�r�^ig4�
6�4�U��d�C���F����%�ѓ ����%e�ͧ����Ҝ�E�'�����P!����.A��������`��ꢺ�I� ��"	�����������cp�g�l$��+R]@~Ǩ�4�D�����m�yOd]�����L���E�a��XlJ�<h�=)�m�,��y�y�<R@�0/Y�����G��6�rR��'��>���`�7�K����E��$t�H頍f--ynl-��_�Ԍn�m��|�ʹO(ɛ�@������U���+�G���Z��Q�h��/�s/����]��JJ��~�mcG��y乶}=��?_�S/S>�{#��ٶދ+((��k?�D��q�G���sR-^�BڮX{��Y�Ssaۂ0'�[�F�_�st�};��%�9��"
�j|n�@������iv�-����$5<����x����7{� ��q�F�r�:�=�x�V���j�V��zZ�]��c���]�H��J��"C��щ���8;�1AV�,�.F���7����!4��I�����e�#"�b��sd�
~zz��J�@8������
��&s��O�yN�P��}��ۛ�}������/�N��,�^S�y�r�����}�ۑ����I3�=��e(�P���O�۬�1W�˗�'�"4/8!�~D�/_���Vde�on�zRl
�dI� f�o�v��؉�V=���G29X��ZG ?`�@�k��.�y����l������E�$�:�����e*Ѫ����_��͆o��U���L��=�������� Vz}�N�ɦWf��	N|�h��N����ݓ���6�¡f�5���ڐ�`mD㻻۫��>�#��Mrs�sp�;$���^+o:kh|܏<w���BDH+��ɫ
�2��ow�s��'���222ttu�41$2$���a�1�K�m��\WJu��>y򤐏���sήx,=U�\�S���u�E-��
Y?��`��mpx�}���������r}�D�*�?}�d�9.7Y�^�=��u)��9�����!�D�k~�������5�q���g�5���H��<�P���I硺03�__ ?Nٌ�֫����?��x[:q_l�/�>��Y���n��gF�M###s(-��bO.�dQ���~uq�W��"x]W7h��T�A>��B,{q�ܹ �>9^"�@�C.b�s���h��r����o}�o���u�s4�bS��N�ss{�����-�哴GE$S�)[&
�!�dm>�F�!0�<ҀN�͛�U�`�s�&�bii�"����*L��c\`�x����j����8�����o����"}}}�3���2_�n�S[�93B,�]�ѷ<��2�_�����H����6� ���S�V�i�p?>y�_�T^����U�"���0N�@s$�?��{�0.Tt��y��Ok�z	�4 U�Tʖ�ɴ���S�:urs�����yJzl�k��C!�̾����9�q�2��Kc^g�
��ȋ��7���s�?�C�=VX��(�� ���/{��m��~��d�'��Ĩ�8ᴴ��+Gg�24⾵Ӷ�0O�||�}��-��)]�v������h2�1`�����F���Ah�|�X��}�wڪ��|��x6�>4����H�Ƽ����@��Y��E�cm�`xz2�}m�̹�ź���S�ϳ�/˯���@����a|΄pg����|ۘ7�ɓoJK��i��K�������0����s%����oIB��=<<�@Bu�G	YA�*�,͆��4]_��h��/�_�Ư��J :5?�@& טY�k7'z��
"���-G?'�9����V��l�L�%��\�04�\XV�,0����w�DXC�XI.�
T`C] �t���ڳ;�]�.�=]��Y
e�	ĒL�I�:)��)l��yG-�����q@��]�����pf����	>v������;/iiM��Ŏ,vi 
���-��+���e�b��/��[P���o���x����B�!b�]���0�Z�p��y���WIۃO��:��	h��O���۬o�Q��(Օ�|Y�}8bW������z�8��@��]�bif�'�xL�N���e;y	R�u�8�����.S�+P�$p�
,�]��A�yIC�(r�f}]�h�,���yL��iCV����AC�ӗ���r���;���i��Ou;�z�\�t��5'��dQ�h��鋃���*Ct��`^���Ni�p\߾{��k�0m�B�ޜ�i��E�\��7o~�����X<��\(�8�xQY~�ԏZ�H�t��3�~��!��r�s�~#����?����%���s�"�.]�Lm��Y�׸�w�a%"�v֗-�(�/6Wy� [1{�����Q����FfA�5?γ�}�6�����d
�Ү���/��Ƹ�ñ�U���A|�G���ɜ>5�|*ÉE��CCC̙99�_�=�s���"g��<ʝ�`K�u3o�i��Խ���Hq4�ˊ_��5������-�黺��U�b�!�v��X�,��i��_O�5׮��^��F���^�oyS��NB	�}��1w����Wo>�.U�o�
�8Sѯ`��[��������-DHSӨ6s�B-R�(D����>H�mSƸ1�܄^XqYKK��6�B��8�?RC��][|/�!�c�d��m�2�$��p��Ȁ��װ�7�~\?_pB�X�d��?�RΪ1F��6�(�F�o(���˺Sy^[\];κhebb�2����Ī-��F�/�c\����;P˅DQ>w�ߧY����_��;#�b	�tz��t��S�ۋ]���oɭ�'Rj�V]�+p������~$9���T�����HR,�*�G�3\d�+~}5G��7���vq���P"gHMK��nd�z$iQ\;8���;+���`�˗�q�.�]h��O%ɲh��w��P	G�ܚ��b��2H�H,ʇ�=42��|O��W1������;y	��L7N/��b��Z��~�����VQ	X��<���v�{�5}�. I�L�B�$�L�#*����7�$���8@�c����)�M@:�5�������|����mʝ���������T�b��a�j��J�-)���@��_�F��7�Y&F���v
���t�)��ĸ��r�)���WL-��- ���{�jy�.�ďX@��\�/~�`�R���f�,K |�[�E� ۟�>H�ծ�����m��$�`: ����X�ȒB��|��^�gϞY��0������jJ���\}T�������(������ҍ	�"�-��e��HJ����t�tw�tw�� ����u��z.�>��޿سgF;��:+�Z�y��~p�7�|i.��~�E��ƿ��qٕo��|r��J*nJ��Iq[;"�{��s�<���*��M������(�@H���D�_�\���	�dk�dv�^G�Z�\؋���:ת�j4F��vMۿ�Yt��K$�ŕ��h���6{�Ĵh�o^��4��1����x�y��&����Ծ�M����⼛�<��δ�+��]�*��7�IF�}.s��4�R�{N̛s� ����`w�+���2%*k��^�ay\�L��:`z&&��$k��8�ͱ����-�~�����{���$N�/_V��8$z˵��,� �X��Nutθ���lw�0:O~n�������n1+?�i9�h��Q=V������B�me�BA��bdxx��p�	d�`ߋข��m�J�~��\�w�q��.jJ��� ��ms��������������<�G�;���QU9t��ݢ����Q�{��$��e���n��w�	�E�\�t�&�p�\��D�Մ����l����8R��j��zC2N�Ć;l�������IH
xV��>S�;���X��d`0j��\v���� ʗ��n�O�n7�LAU��x:k�����i��Re�ot�.�L��B��@�:Q��b��q���CKn\�=�Ac�D	+�v9���4��l
x�U�Vט�$a����t���5	
x_���ǉ6�Mf�Ӵ���3������ߺuKp�"R;g��1
;�i�8�Դ�����a:��`�Y��og_����65��eo�y&���BJJ��$�ኇc�jF|k�a�ϐ��8���3��rW;ށ"H�Ծ#�A����u�E�;w�|��3ߧN���o��	�4lڵ\�	�OL<��U�E)I:ن?������,8HKK{[���!GѡX���љ1j�\�����@���m�q�n��л�Y?Ֆ��:��o��)>YPHH���fB�CK�8���Б����ˆ%=��I�^�X�h>�t������m�lm-�7�J���yo���u&�o����M�y�������<���<.p�5�ß̢��Wf�y��`�ǐo�m`9�p.������D�@��-R���ֈ{H\��إ�Lw4�\�-��d�[ԩ���.5��J�aH!�`_�ĩ�|m�S�r�I�,!!!a���j�O�!�7��kZ�Զ���'Vu��f+�c�
��I�� �ށd�U���z���g#��=�!
Yz؜Scgc�7,l��2[�+~j�!�7JP�m�uc@�!p�z�!���\h���%{f�QT��a۠g�efզ�ׯ_z)�{6�x�,0���BB:w�+��G�����o��h�sj%:R=��M:-�VQ���v�T�-�u���t��A�����ϣ�[z�W�^L�;��w; $n�f\RT��#��',��|q*P�`dQ�r�~WTh�:Ȧ� ��`����a����ʘ�����57b�¬Q�R�t"
5��� B�y�۵�* pr�)�AH�r��s�#:�����t�VdED<E����8����u�vC�̍ݽ$і%]��q$frz�C[Ձ8��E8����ѽ��
Ix��:��O�SĽ-�"�:=�@+����>z$K����z�sT�P�=����?����7���)�W���q��l�3����iii�jeG�<yr�c�=�������د��*S�y�?]Ȼ�e�1ӛ+�Un�؍e���~�~��u�>#1 �ʆ�t��i���qٟ��������}ͳ'$$d,�q7��hD�!|9������&�+���E[�v+Mj_!"�G��G�n���p	k�jk[�0[��#_�J/h*�{t�g�6�M^^��b_n�;J�[$��*= �u,�쯞=^�*j�XH��l��{�E��lV��>K��JX�6�Iq��R���{!@j���dh�y�`�yk�l��-��9G'�q�M��J &y��*q����E9�xI]]ݗS�	���i��850���G}�Ap������Y��k�/�WCX|�=�_�}�"
���,�����y�}~]��,53ߩt}{�<3�Y Ƴ��#t��A���,)t���AG]mlX���û0��t݁y�h�^>��Jy빔��`ɯ3���馦�PYIt� J̏?*�N�s˂%�f;��A�k���Quuu�dBCty����'wsU@� 2d�=x��_g����!W
!�����"���E������X������o/RǨ>ܕ����n��AA4篋�E�@H��χ�E�-�^ۯ���m�o��[.�D������b�f}0Ͽy�w����1�	��S�o��λzno�R.@Sz��K'$$|�
��.[<+���i6^�戳�	K��� xI]`-tuE�#/���J�3r���n�X��"��kSr{��I�ݲh���S/A�.�0�8t�Z�h҂�\�ל�@ ���+�;����>�����
�}�Ǐ�+ʋ|�Wj���B'm1��f�Ny��ո�̕YT�k1Ĳ�AZ�Ha�XrN�/�ς���~��_e�Ҁ8���j$58N���53��Nh��S-�󂘴���sA�z<j�/K�¸i ��ꏇ@���D��� �4�i�����1�����

����� b	�7������5TM�.��e_�+әλ���An�577w����=|���OBs�� �Y���\ϐ5�c�&��#.ct�7�����a��=P�g�cw�:Å�������lb�����!RQ�����;��Z�O1f��F@�e���ht��ۣ��;����~�������"�Y�s����Em9A�S1r��j!2%<�H#�&@L�I<<�6����U[���5����s��F��C����;���(��9����c�>ѡ�%@f�;��k0��!!YLe�'ͫ;�ԩ�wsS$:�܏n������m,dgg��*�Hp��(�I�'y�k+�-�u�fO)���\[��w�6x���N)w�=�.1���ʿ�O��>����o',i�[
(�DWo�r���]�hw���������]$"��}���˭���k=j�t'�v߻rE��'�k�Ĝ9gǖ]щn�{Z��{�x��BŴ�M�^{���׃hG�$�_��|���f��>�����ü�h�� ��X ��=��y�����O�8�@�&�bu����с�>S#�����n�S���A,ӫ��h�E�\�&��S �k���-�a�
ہ�{�W���a�|�S�F G!n�t��.?Rt�����|�F���O�hg|��������eof�wJ��s��[�A��6-���R�Ac��T�k�~j�S00H�� ����"�,��{ ��ƅ������ix��? ���3Eװ��.s<�Ob����Ak�j7�Q4q���8]��|��5�r[/� f��P���� �U�V}B� ^�KRV�����Bz�P	�MF�3�����������>i99!mqQQ/��7��r��[���o[�4Q���d`�-�w_Yo���JУ֨	���`��M�<V>�L��
���'��r!�:~�������ԡ��&:�� 5���˪���-��������������L�x�y������pϝ������G�zċ-��w����^]]]���������Τ�����L�����/0��4��E��\�KU�"?��浪0Z�i��p��
)E[S߿�b��L��=F?n��{�G�K��Ʒ�Ӎ�z#�Ή��.�	1��Q��G���?��R7�|)�A&����h@#�9��+��ཛྷ�Lѝ�_b�*Ĩ�&^<�],���\�vG�R��"��9glL��vQ���&?I���$��AL�7���C�+���R΀�����Ni{�B�z��5�.۬���v������#�i80��m�UQt���Ǐ��N��"t���)H���&ZH�%S>�+�G�w��w�T�����\��ߴ+�y<�$D *�s�2l���^9�����"3���>0+�`C"!$��j�����K>t9��s��Bب+S��qH�B�^���c3��ݑ���2S"�#�߳������@�4�c�����?��R��O.�NK�"��jJ�u66���atAAA��*f��� ~c����yÍ�ˇ:U/�?64LQ|�&E`�0:ח�V;�I��deeU�^����)�6��:u�����^�N�PάA�����5��+� 1+]N�f29���ﮃv�����f�E�*R�������uI�@�޳�4��{IЉ��|�)����C�
���6.]��)i#
�K����R\b��J�S#R��O<-H);Kߞ��lqQ�)�4�S6.�etر��"6��_�t^�Y�m��C��ڬ�H ��9�4�R?���
�,�#�?�w�'ɺ��6�oN)���_�>�؁Z���_v�o�Y����c2]Ml�;�G�C-�Σv�m#��gd�W����O�x�����`�7)*7K�x�]|��L�l	�������,�b�LxCP)��>ˑj3����썩���NQ��O����(�S7M��B��;��~W����бj�!�R8ۥY��$�x���N9 G����ɣo���R��,N�5qX�P�����V鵙N>�B����4`˼�O!���SG5�-u�e	�[q��cЯ]���o�y������(�(��}��2������\�rV��jA�������C�����;�;�,Cn����8���ħ7�,��ׯ��?�#ɸ,*])��6M+�=��Wz��:����V2���xgP[Mm(��ε��}�����1,�g7	}!����? C����#��ͱ�$9�����U��C��E��Ԓ�����&����������Ι�����⵻�.��9�0G���&N����[��堗գ����M�������SE]�H�e*k�~ ]qz��r�]�V��gE��NO�����܇---|	))ʨ��63D��{n#$T�866f��u�r�:^���ޣ$����8YV�YVl�|
�,���ۯH$|�:�(�Zw������8<>�Tw��5���C�H��p��q�NGW������h�[�9�^h�ziwޑ/j�r�ұZ��7����=k��j �ޣ��) �kڿ��F�d�~~��J*4�М������*v��=�^|�2ǰ��I��L$p���!�g�О6@֏T�n5�$ǼH٪�ɸ2�(��wdԯ�{����8K,�NuvʎG�;W��'D+�Ͱ��l]�Ұ?�Af#NX8�O��5N�ڕ�l��8�#�������7O�S覀^3��{���O�6m�Y��N-��`F�������G�k�Zr��s`�A��rZ��O�O�tɷ�/F��W.��[[6AlFa�3���q�0|9u+���-Z(����r��6q���Va!��޳�O��m�|a7�4qħ�f����.>�TM�7��mȸW3��(�O���QI.&>^/~5��[��I���!{����I�E����5���QɃ�qog(`��U,	�W��jѻ���+��g�-f�ϓ7�>������n�h'���oO�����䪕��F�xl�*=I����й����0��>�l��6�j7�RAW�"V��
��Bvz��J3jAgBXL7qx��MJɻ%"u8�Ef������b��UI�(�Ɠ/bZ�9@T�.�<�}�����;��q:�,����/�|�!�h�����T��=R���Vٔ��.�m
�������9���O�tA|�����Y��l�2k7����˹�;���j�W��Y���Td�\o�^���t���Sj�[�X����CF��3�Fd�f�/Kș��S��&>g�tw��؝�,4�uꗑ���d:��a�D���| L����;4YE&��l���P������č�����SV�����~]2V�C�r����UaḶ��5ytS�v�3s%L�o.�u�s�HI��}��jЍ_Ihm}nj���Q�X(��Yrن��K }}}���eV��ܯ�u���w�{y�����^�ǻu��������;�m6~ݺ	)�|U�{p۽�Ұ������"�;��^9�}�ȹ�/�E5�(���0�7��M�rN�1<�2��7�t��C��]2\��D�� �4��_�-{w"���ދ�?k�!�����A--��Dk��w��0��9�抇q˩��e7��6��u�n�h�hˁ��0rX&mko[>ߒ0�/iz���/�Pqص��	�n����ffC�f�'' &R,��
����z̴e�q	\;5�F��\���'��;�������R���\���3�Qߔ0f����)�/Gv�5�b�~���1r�+��/�D��X��m�gӨ�!V4.����.�ё���Ϸ��o�t��%N4c�[5�>u鎪��̕�_n�����C3�<k�e[��� '��m���{fJ����r��ŶbjGR�d��۷�ֺ0����9�ž|uqq1�_Ev(k������d���z��gބ��T�����!�����t�|(���;���b�ݣ�����*P+��%#/��Ub�3-z��v
1�Ą��d����8�~�� I��~����fm�������[|ލ= ����w��J����M^���w��Lr_��H�TT�oN��/����5��S��ᆯ��bk����1k�_V�����֨��C����������pǢ���^*Jʕ�����\�TЃ1�5C�ܙF�@��߶m�����54b�[Z�Z�X��_����1,��T�|ߒ�w8�>�����P�5aA��[#�A��OnUV>Aߝ7Қ$��q�L��?
ZfY�S�i���w�1'���N _��<6;� �&��#�Fd J�Wc?����gϚ��K�|�����!@�s�t�v2���.�$�C$�!XJTB�{Q�F�AH\\FW7�@���t��YO��u�9ԑ�g>�bZ�&���H�|Vu{.f��Aw�f!�E�(��L�����{G��e��S^M�W�Z�x�x���6k�7ANDDD9)&��BI�A�m!i��"������YL���ѣ	t�L��7��[׮�4�B[��8?�x�[��c�`����lr�(�����ժ�*�(oR6C5]]��"� ~R!l�4�����2��4��@/��U��M��cp�q��=�K���	{��=�x��А��=3E���m�/�0&Bs��Y-�c���T�z�mv=t�b�\�&��K�d+>w����01V��Fw'#y�DP4��#�������Ы23��L
�q�B�2�F�zNv=���TW��Kȭ�M3p������{�9�/�Ys�'�+*�Eg�����^ZZ"�t)��ڜ0@���o�V��#��n��G��c7�hk��%��N�u���X� �e�>@����0LE��Z����w]ؘ9������|Q�L�18�}U�c�|�ɴ
r�6#lz���LLL�v�zBXƟWكԻm�9bw`_JD�3�I�f��z�-2˴���śuF�,Z���.1�t��7�C�ߔ�y��7"��_t~��֗��wúg�@W�ʤ��R �+�W<6::�>�aT�3�`6Pd��1�:۳����߼��)��>o�ru�O�Ag�&f
"�a��S11�0��8I;�MLL4¿�}s�΢�<Ŕme��,��\c�9��d��Vܼ�E�z�A��iih��Hz0�V�U �ꬁ8�A7+7y0i?d�ܙ���]7kmm��m�����]�Ŷ=�+41�7�ͥ�	*A�)�qv���}ċ�}`��ϟ;s����{d� ;�~�Cv�Q����t�-۰/mi�4�V.+H�U�jȹ������VJN.hƘ}���|���>'�#_{}�o��\�r�EN��^%k�g躼��d��y˙N� e�������x�Be@�Ǐ�H�J�&o����[zO�m"x�le��lD���C|?��>K6�ثvsq!����e�e���f:?�nB�		K��$�`t�kF*4�M��"�h+�#�?��4����F@�0�d|�fuc�G��.�U�(9���t#V��'�>]�ll2 �<�1G�Q�b���_�t�c��1�\v�o/R�����R`*��nT�P��t-'0�kO���� 9��|��ed��o��F�;8VVUјC�(f�����KjT �:����b�	��|cA�EB����vڗ/�YXYu+?\��BS���O�����o�J�Z�l,��L���n�v� �<߿�f�zu����X�&�#$:�0��&�C�y`�Cxh�]{�.�"�썌��Nڌ�Db�k��O�?��!����A�q=��{��3���5��!��q2���4������RQIE=d��uG����1] %M�����qX��=V�������v���5�մ92]����Acv��1Ϡ�n��ppp��*�+�����a�v��,T����Ң`
�=��M&��<~߇�ݙ:ѣ�/!�{�3��$%?��wF ���R��s�+y�L��8�Ç�-&;B=�T���|�>�5�"?�GE;S�ײ�&� �>w�\���Ͼ���ݱ��5c �8{_c�����Wۦ#7-M
m�ە,�be����Ĩ���m���ʇ*��$+:�c��S�j�M�zF�VK��Yn�����pf!Ǯ�	��}�j�l>�Х|�QR�'V�0�������{�2!�}҅������w�8/��$^��	 ��b��3���tz�cJ��������]޽�Y�h�e	�h<}�N����H��3�� ����i98���^�o.�h��Iz._�EC؋S�N(�i�~����w�����J� ��ö�?�������BN�S�)��y�A��{�| Jm�>����B���0�q��c�?F7=h�k���#�T���
V������X��F�ߞlj��;@�r��=������Q_Skk�+����~��emN��|��i�� ��"/�&-mH.�\G<��ȟ?��@[qqq9�"�)��Mg���D�nMRդK�k������H��|��vD{vz�﹖�mY�7�z F�X[��䙚�β��?P/͉��g���!!��=/�R��W%ϕS�g5�����\��W��5=���6.��yz�]�O�����p��33�,
v�t�r2���O7�����)`h��wb�SOOb�|�̳=��~�.�vc������ɛ�,�k��Z�b6>��E�Ƀ�A:��^�b�5�e������w���zv ��7��oM��z#`B�GrP���b����q������.r��Bc��������-8C��B�Py�.?|P޻w�<�Vނ���;,n��4uk�'0	0�7oݪ�n�'!#��b.%���y	w�nA���+�{z2�U�����������_��g]�p!����~��p�4!!�+n�=M�ByԘ���߿��!�S��f�"�6C�.���aQ��?��4�.f���Jy���ge��Y>��z��&�A���8�{��'ǨÛ�K�3�
#�ۇ"�C�V�i�Ȇ3|�����]�~�C��#��Ds���jH�v >�@Ȣ�NbR����ײ����#����y�S;B �o�$i��<|�0�a�K���
#o��f�9�q]�.��֯���r��(���l��y�Z�s9���鎤����nolK8v~ ��u���lq#G<��f�t��=|HJJJ�z�A_MC��� v4��#ᵳ�65]"_b���1羱�a_?Uօ�AjT_��j�Y�'�YS .��Y3���c��%ӫ�]��~h]\CC�����"e}Nl�4<��|���hrz�<i�gV+;�r�0�7�o!b��k���rN�S���˫�:@1J�>��� ��[���Z�����!�9�^ �[uz����ڜ3T�q]+����Jt�e�S,6u/Ş�L�gߔ�����{e�������	�8q��wϱ7B�#�O��J��TTԫ��\9� r���c܂��
�:-S`������:�ۋЊ�>kh�9O���G?�@��y�O���Hv&���E6/�n*O��e���T�����$$	:-qHM�a�KJ��W��&x
�����9a����-&��S����� ��Q ��j������E�����?J�hl�����],�?Ɏu�����`�BS��t!(���4~GW#�kR>��.�.��0@p+>���B��&�$������o/Q�}��\bųdd}�1Ԥ�����2�y2E;�'��u�̫��������ׇ~���߂]n����"nk±��o�����i�~������˫�ys��\�]u�����'�)[[[�a��R�f�^?�]񽲲��?���2� 8�C���_C>q%(L���t�{���{�@rq]�`0�
- j�>�`��;�L�3��G�\�o�#�ᅡr�=�^V�Kѵj��e4�kЕ���Y:��]�;1!A�h�	�4x�6`~��$�t[k��[�n=���a�5����">��@ [lL�e��r�X�-֍��FθFצ{�S!It��3"22�l�
�<���x���������8o����i/@V��5S��6BS���C��8/��������*CT���z�=/��Bۜ��tY�Iכ?��񩈆�N��� ���������ӊ�`��J�(�(�MP���q>|�t]}�ܤXBW7���o?~l��ի)���!/�Ӱ��r2�������Ѓp���v�!�0}�P�En=J��G4�Y���ν���gZ��+(�����Y���B�9�x��H��j�H~No�xI$��}ȓ��	�>��\�����"R22�SI�{>�L���� e��̷�VWW�K=}���-���D$D?�r!�W���Sc��)\R����	����aL^�N�{'�o꽍�v|��T�-&��m�ޑ��!���o-�F�E���0���"��"{[�$4��;��&��j�3����Eb����J+ڗr�@�f�z� ���qT��_�~m����M�_q�Vx�\AFF���E�ǥK��0���������0�2Yk?��q�'h��#=@�Ƥ��6�..�� �����"E�����8&#5r�Q��u`��M����L�q��-�������-S;W��P�l+���f�c�7�����5#�|��q0��@p�{k96���/����@�X/�x��<��1��/_���vA^bտ���#㳿H��=�ʞ*�&椭��+%Ĝ�����k	��/M #�ܞ�|SV^�3000�@}{�3�+�4N����77���}��ԋ�~k�Zգ���˗/3�8������Qw|N?H�����BCA0�9t5zr�ӫ�B��C�M8C��\�v�l���)�G�@����i���j���j~��~���-)��}�vE�[�>��.�Jw~8��i�wH�@o��-����x�Wܰ㔁�!�sș�s�t;�+In3qU,�$�K�8Pl�+ݎ��I�d~+� �g�8�; @�&P��E>� �����X��Zn��3����B�
J���������QQ @�II}��#��{"(�U���R��]�c78.{K>�8.���177wk���認� ����_�%��?l�i��>���\��11?��1�F���"ǵ�-�Y�J-��	�8edA�rJ�NQf?$����7���t9�81=������y�vj�W�<#�ٵ*	10ys��֮�&���;{y��aAhv�潧f�}�h'�\�`.����(�r݌�ׯ��0*�R�>��'�ĵ���n�La���d��Cs��7sB��;��e�ߥ*���y�����U�X�);�~�|���Ғ��Y���c=�:�
��>�[t�qq��`��+z��]tF+?
	g\%�l���{r�=�������u��Ew��}�0w�����]�U�)E�T��6���M�}=Z���#z{C�M�bM�����z#do_�3Z�'��Mƣe���h��]NK**~�d��9��d���Nm|>�O����Z�}�ϋsG*�[$����/�Yf�Tm�!�� $&�6��S9�縿��0�	�+E6���\���4u�,���l-�PN��#����zH ��E^f=�d�MÙ�쪜'�6�:G���ʏV�b��P�g�NA vrȕ"[��������3{���-@��ڄ�_/���Q�n��&>9�,hwq�C�X��G^^&��ꊪ��̌~�\���-F��-�E>*ݓ���ʨ�g�
`cW�?#�zYS���@o�`���{y_���?�(��{�Z[Ay<9����5o؝V��USSSUg5*�c0�k�x`�۾������k�|9v>Þ�n��N��N�ᱼ�<:���+`�� ��p��^��y�N:٬>�+�g��&=�q�~�w�s%$U���\��=F�}���܋��!Ă�V���$�W����8���rj��^��(@����K#���g�\�OmPX�1�\���S�K��F3 �	 ]iJ�
,�ҷǲ���X��a�H�i w�Gj��X��?�q�Nbjjس�ϟ��<�a2��>M��\PP�.�-M] )��x�$�ޯt:� o,?�V������n�^ݓ�1�c֨&<ik�-���6k�->��,:}/��g�br�N��f��SBv��ڭhE�/�R��;��kU�Uu��[9x�<�:�{?��i��t��%��94Ԁ�?��`��WEE�7�w��l�Ll� ���n>�Y�*z]+a��3�ߚ����c!�e��?�7�.Ow�jxP.y_�B�+%�%�ה1Tz��6�g>�o7���%�~ۂ�3������Q{w�|����=��7�6ߣo�XT?��I3�N��_>1h�d��6�~{-N�Je���fՑ��F��gIIkԹ��3���Ï�oMU�2q�E�� A����C�T9��xS�$+�$&&V�vz��%���I����B�ZgT��Xs�	���%�5ҡ:1|�Z�kyd|�M�Z'a|�i�|�d��ǎ�,�����_o���6̲|��d���W�Fo��
'ɤ�������c
&0((AIuM�'�	m�����zteh%!�ya�Pz� �T1�U�P��� 
h6g�p[�0�nפ������ʤ<71I�dw�����3-X��O��.��^�L��*�%O �7��S��Z�TT�8�8]
�&a��d���1l9(��8��c9�@�袓�v�R~��	x=��l�z ��"�c��ɜ���M�k�!W]_�τ��-&��t:a�b����W��l�9� R������i��D�e��.�]ڒ�5���JBLb�W�t8�it�����i/�O�<	O`����SZ�oOS�jɎ�vzõ�.�D1�]���)H�Ʃ�$�W|����@0e�r<6+�?LF��� ��ԝ�t%Ԙl6�c�Gh�akڑOyy��r��~5c�yߕ�OUIE����v�˙W��IC��6M5��j�W���0+<|�f��q�! :̋65�|�9Ş?�S2��C44�1zP*���}�'w�/مl���L4^E�kk_�x�@R�����c_�o4�|�^)�@BZ�
ô����*�ʀ�oIר��N/��+Y1��I���d+�?hq�nFdȚc��X��]_0�zXK*q��&���~���������� 8@`��6���G��1��\JJgw���#��zY�=Й��y�fa��pH��ˮk��~04���qT�t|�!=���>g���`���^֫iiT��u�6�1vu�Q�5����3�F��Q[%R��6~	������/O��] �^��x�+$$��МX�����G�s�"AR`2�O�av�$���]L�/ׅu�(qq\>���W�7�Z��Ł9��>4	ld���#n���ʅ�UUUy;K5`i48�-x�021I=}Z����]Ů�b��䋒��/t�;M^�Qkk�M..������3N�={qө��2J��2��߽��Z�DKv��/rb0�D�TX��/��ho�����]��oI`5������|�3�E��	i�݂��0�r�KKKϟ>�Xn�S	P� yl��Υ���]���:d�9����`�@(C��UZ��c8��u��в��ra��>j�F��U��V?�w���V˅������Қ���޽�]{�ϲ��B�@P�hjv�+`���abZ]/���)��k�Lj�z'!;[����
M6��㨟Z���eO���o0%]�h�a�� ������ˁ��߇Y���&k���01�d��Td���7<�����`jz�sP�u�vm(��|�|�G�M��ƨ9�<ev�I|���ɖ1��3���eee"''�ە.����v�^*)�H�>��y��u���ۊC��y6�{3{8��������æ׿K�z��$&��,ۿc��U߶,��7�@*��{YĄ�F,�bϟ���9��#oa&`H�
��%!��3&��"iL����q�����r-���X�P�B �e(����@�"ۮBW���Ft�m� ;�P����u����
����kq����:��B�:�=#���u9��L9C�%�¸h̽�,]�q�ӧ�n�>��8�Y ���ѯwS-�>�##��n���/��.ށ?�M���t��]@Ω��t��nwƀLF���'Y�C�Fv��c��B�qw5o�^0-x{t/�zo��������]2��0�x(AQg=z���D"'��U�ڈ7o���]�j4P�>���I�3�I��o�
8#Zq���QyO9�]���"ϝ;g���8A���r�N;�A�8l��(6ha����$���L6��(Յ��+��J�߱P`�����zcނ̧��S"�`S�i<�D�?�nF@D��Ny8���nMw�~[����T��:�"P�9:��ϟ���f��GN�݉�復����iK�a@����h(�[=_��  '�`)�32V�w�����)�.n��o��;"�a<���72c"��+���0l�?�M�)C�m�ey��M��W����s��l)R�h���컛?�o¨�r�'��˫L�luU�&�1++���AFL�LO7V���xC8�V a�?YF�h- ���J�x�B�\�jN�^G5�]է�7��1%]������h�ې������D�Ċx�?�}��1.:ҹ��mr���������~xX�Е���D�TeT�洜���se�"�����?��w�N-*RF�6����H�G��T>���0�� J��1�7aJ����j�1@����o��^��+A>
����L2��f]��u��3�"�1T�x@[���F�c�9AdL�5�7��>a���+*~{{
�_WW���f9�����k�lv���,�&J�X�@Z�k]Zq�%w���IT���CK��:# ���IO��U��xbR�����3��˧JpG���[l�8Xc�oG�&9�b��5�1}ή�����>�<�Yz2�I�U��W��'�6t���0���@ ;�2�)7d��m���qbع�Z�nB��j�-�>2����kws	�孪�%����5��������|2'RRR`��vFo�I����zp��o.��~��ll�]�X|ލ{��Qwƛ'��#�)�%@�f�GF��_�4%�%��T	`��k *���k�&��v��?�TAGq?�)\r]�݇�ld�;Ñ�^qT%��\]���r���uoN��� ��{5�����aff�2�	�,��9����=:�c��`F���7�Ο��ucêeQ�BM�se唲���
�5��q1Xz5���eq�(������X�V����;�T6�����[PI)i�ͱ �CS��o���cΐqVzw�~��) �;}��q)V��◢��1���h�X�<AEӡw��Qu\����E�h�S��>�v���{E-*ƨ��L�	�;��N^Ĝ}�`<���>0IУsh-F}�R���ETt���)N��[44�A��[9ur�8'��*	11�TVl`a9�Bњp^�>�:�#����g�0����g0vI���24�g�2D�0ᨵu���y*~�ƥ10~ �a�4��G;��8J\x�O+R�� ��@tc朧�O]��@:ԉ�M�s)Z"c��?�&�! �pqq}c���Z4�abQ5�֭j�'|&SX)�`�1@�>+�ژ�)�=�o������-�������g�+� ����jo+�c���N����$x^ggg`1�k�'j5�)c�[U�ٖ���V� �|}���������|(hT�rŧ���]X0F	o�`"��1ȋ�"S
^^^hi&-WW��X��8��St��8<��NwZ�!B��i���s��(��s[�#����,���򟺖`=�'�3���R>k�s�� .���HFu�56`2�@ZN 0��Ł.���U���L�h�� 1�� 6�����sNE6Q�ϞEA跄��J��{�⅘�#�nH@@p��#_M��i.��2����T62m�p�pG�W,�"��o�k|���!$*������+.���\\t	�κ�~�%	���M<��f26����rˬ/�UKk�$Rp�>�D�k�x
ђ�����ߤF�d8�����p�-������MV�5�bN�-�q�(�yM9������q%����K���-��J�6��*���ƶ������!��$$	nn�Q�t�g��v��l�с�ί����W �ӧO�/J������y�v��lbR�A�4:�K�j�x�A� q�
���^b��;@r��8����!R��0CΓ;N�C������P�����|!�4x������ory��9t6�޽{7��c�������0ڝ���	C�%�����?q�C����m��"�{ ����;
٥�}s-J�F��(AÁ�I[���Z�A)�  2�	{RdLՐq�y�ÕS�On����א��g�^�]��o�?���D�xX��㶂�@�VC���g��-���5t���g�ug�s��tj�|��1�*��)�
t̓�o6'İN ��3֌�r��B���_�0�wqXxKq��ݴ.3��O�]9��|dq����?���w4���Vl��؄̂���^�N��2oֲ�3�R0݅ͮ__��g�.���3Ja))�F������m]�S�q�-�Q?��G���elV&���A����l�:%C��TR� �aԨ&D�n~
Êd@Q���i7^�]�q�K�,��4��˟�� ��w�#;�~����T@>HP&��ER�a�b-*�[JZ����w�cu�顰?]Zro�A+�D#���l�@�V��&�Q�_T5����l�D����?��dE4LZ�~-U
�EL�%u�8ήv����lيs,�^�X��ฝ���1��(ir{j���?]O �o�n��*���`ǀ�p~�E�%xY�:�I������!��WHE�d�H�����+�����Ә0�=����[7�T�N�Κ-j�^M���F��b�z���V��xD��*X� `b3���у�s<������!���0r�&��2��7P^ݜ��ՠ�Ê����R�ʜ�.��N�}�� ��6E���@g�� ��5HK؋��0�X����9�N�Y��RG����i;�z�����X�'	Ө��9����Bt��3� �!!X�6�{4��9�}��t`H���ف�be�U��#oy�:m4<��z4��g��,��į7���vr�/8�`�Ss�מz}:%���B��)Z`��k����ڵGfj�����Eh�����X_�4�A��+�jos|����da>��B�b͸�����4+�Aa��M�nf����jw��kt2<j7��7V�^RC[XXc�gj�®6]�Zf�l���	�f�l�t���ק���K^���C�����՞Z@j���N� �����r���Lj����7�x~��F0�_4����'�Р�<}���G���FI���o�`k}�h[S�c4�(F0�͈��4)@�A�o����Cmq�A�4�S�a��|�.ƶ�v��ƃ�`<�����Rr�����if �[���ؘxЍz3�i���y�I�B��,S�u��wh?��f=�:��*v444�Gm����M���;j��X^M=wvqٺ���ݽy��/��ж�3'2�p }֫����)���1���܀�)���8�~��
����(�>������0�п<���+�Y��M�.T���ؗco!"≚��&��.�-��H�fGߞ��!J�u�i3 ��.�OeUe_c{&��F�wv�)��� �x�ʬ��x�zD��P��_�Iw����`o,��z��uT�E����jPoss3�I�[\3�[׮��c�%/f`kg�!d�[}��5Z���=��
ρZ���ͨ#�5���K��E�?�8�c�U�z)��/��Y�� .��kj�,��tt�U�{0��Ǎ���SiG���R�BN��***� ��w�n,cm���g�1s8m�o=>������dd��hCOp�\�Q|�O���"ݎ����f��Y̕����ޕ�5u-�[��U�Z�,`@AD��,�(hĲ��QE	�@���J�u�TR�%��U��f �[��%�@ț�������{���'ܐ9��9���f�̙�G�j�`���>u���#���˗Q��כt����|
�0B����d��� �{3:z�x����p�`w���B�aFF�m/u��Q�L2�n٩ �ş/T1|��� �!�R?r�05�Bn��F#���0Y�d��g��9��,Y�X���.�T4ڲ��rL۶��eVnIE�������1l�ʓ;}}C����a�v�.hَ�R��p�o��A��;r-�Kzp"^�Ԛ�1��UGk�:��Uj ���U,(��
�P9˩���ASOo
a�/QGk�v����h&���4j���r�.n\=9�ȫ1�u�q�+ 	��D����>0׀.A���W� �Tu?)	e���,/�F��09��
l1��>�����*�m��P��T�EaR��b���'����;����؍�(g.��'ǗO�k��	�5""�.*��	�S2Aɣ�Z � �I�S�Ĭ,ë�7P�.�z�y�X�J�;p�DRǚ�����Tj����%��m���d9�0b`���K������H	�(m{��+���a
"�6�7@�V0p�]w�J:x$�s;�����^;1L��b@���z_0&���=S\�T���`�+��~}i]ޞ`og�����w�yS��?�(��?�������O,��ٓ��\q�ZzNsN$�ơ�n��>��6��lcS@؅�ya��'WU7��;�"��XH��&!!��%h�$(tr!-��ח���b0�R���6��V*h<d�����M���q�el��R8k�����S��ibt,�I����vD[`n˹�7� ��A,�8���x{��`�?��o|d�S,�IիJ��s4i�K�MiPY���u��[���5�̞w������������e=�^A����{���,��\eu�xP�nU\�EFFF8�� �C����i�9�՗_&t�cu�I���B�Oo�XS�_�9��'���!��B��ҭ�we�"Y��U	
<*�R�R����ƺB���OiS))hЩ�F-�}���tk�g�d���~����ǌiow�A"��~LEE�����&��dQϪ��<@8�ɻ{`D����Z�5���Yb.��(�u�nғ	y�P4�Qkk���\Lv^FY�h���g�A��}����n(�i25	�c�Fj ��"�8��"o�@�k�6�ڼ���O��o���N(^��12Ŧ�}1 ��-#k*1
���3�=8Ҟ6�.B1/����L*\��&����?^�R�lHƚ���^G��#%֥�z���>;�V�o�y�ui��$����Q呾2�MA#T�ڧ��Т�k�?���_?~���g�Ș�\�����m�2�;�	��P���K��IjlJ1A�som^�9�5ľ���k����@��Mks�����y Hd�~��4���QzM��K���c�>jn�: 9�<���we%tq����Ͼ��+ 6w�G{x�oJaJU����Nk��D(��Y;��jc���[���I���\jA�X�=j���w�;�|�����t ��;	�4��1�o�U������q)��[\aEY�G7S�-^��<�0l{ɳŅX�V13�C^�<&��w��Uk`�0���~E;�"��F��><�������<~,�s �3Op=����b_V�.5v�f�vRo^[<�itHd�/���*�_�e�h�YE�6Q\�|�^I�R�ֽ��3ؠ�>]�
`.�W}1N�٨��;�4tg�"�1�;�z���e��{����P$V_?GBA;��Դ����=�z��k���*�~�m��e:5�t���O>L��upw*Ʈ�WB�����$4	pm\�լ�^#ŗ��f�)��f���S�(�M.���Ӡ�߉�[Z�r�xG�w���;���3O�i�Y�����K��]��u�w�Y�7�c�#��r�X]v�!����C�w�h� WdS�4���A�-��`T�';:J>�W������m�A%�^|@ި�n�g_����fNY��^�-�xy
ѧ�$��Rmm=�z���� ��Ͻ����T��p�d�&��B�S�W�D�B����0�Ca����0x�SG����О�E[�6P���ѩC������ S�=��`��-X��`_[(���m���
˹\{N�7����4.�[g����/�1D�z��ؙ���9�u,n���m0��������8o ��K:k�7?}�i���2��?Er�V����wT`���B�����62pR�\$;��į�����i4ư��"��A��|��ja3�ܸ�y��,��8�Lv�͍d^��RQ��T&��zL+t�Q5|����o�ս�8!��m���̉���۫������qd3^�=5��;M���o����8�3���ߙ#�x����J�ĩ
��#����]�^򧕵&��n�ΙN�a�z��Y.�rb`آm� aC=>2_�rc�G:��w�"URω��*�I�@J6|@1L��b#��Þ�O��Š��Rf<#���`6��"�ӕԷd�+�$���èQ0V����|ڤB\��V��
f?+p��v����/�8=w�n��"��]��B��!®�d#�`:�+-e��FZ&��`v��6W||����)��@��EVJ5�R����x�ӂ\{Ir�i��ɓ/�G��0�4��7���l���ޗ\���8NNN�n�v��Zo���N|�3g<�N3XWu����γB�cVff�����K�>��ǚ�%����>-�osQN('��	�rB9��PN('��	�rB9�H8X�y�|��6���go�)�����ˣ����w�p�2�љ�����>�7�M���B������?0���C3Ev�u��f���r�@o���A=�$hd���E����������f���]�t�����ak������PK   '6X��g� 
  �	  /   images/4f5a6b59-a216-44d1-a198-112719b334c8.png�	��PNG

   IHDR   d      X�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  	�IDATx��ZkLTG�e���	>*���M����ZMl����iҪi��j[�?jb�c���X�hml��1��b�A� � >A�
"�"����;8ܽ�h�Bz�q�;��>gf��^�'OV�a�i�b�}v�?^���W*���{`�
� X/��У
���			���Ǣ��M<y�DX,���,����v�_�GL�����1bĈ���^o�~εZ����E�l6QQQ!z��B/^,���E^^�=&&&J���������GDD�N�0��# ��[�n�:�N{0E]A|		�� ������q�ƉK�.��[\\�p8�Ff=�x��SSS#��;��YWW��1YYY<x��������@pa�$�LNNv��+�j��@��ӧO[\\�i����;`Ȑ!b���F%y4�KyR�w����o�����;�P����ݻ-Z�r��=QYY)`���ŋ�B<�����3��*CQ7>kt���h�th	�������?��ӧHt�L�"�mxx��q�m�����ߢ���j�9sf��icK�ǎ+8)����F�������?��;�-[v>77W�����g�v�x��EQQѠ����z�J�ǐ������p"��9)�����_]�3fH�_�~�سgϚ�S���>�:- 'pɒ%�\�Rg�J����H��FFFF+A�0���о�}���ȑ#A�c�E�����R�|&p�ђ
�v�L�e�������e����Ž
�ɓ'e�6���
,%%��~�/_6ݏ
���G�n������נ�"?�a�>�
C�������bt�*�c�C.�4i�E���[�|��իEII�d�رc�.�gY�n�'??�* �[�?^�ť5�(,c?��J���@�j6��k(�ܹs�J���ƍ�ki8����T�Uz �WUU%EEE}a��O��@�|�TߩT��Uׇ�"�Z\q�ڵo�o߾�-[�t3
��v�F�+�����ͻ�=�hGAa���U�V�6O��P@����/[
�B�(D�S�T�}�'��;��m֬Y<�6�fϞ������>x>��#�tX��v��h�� ��s�Q)��y�w׮]�G�޽{��_UY*ĐP�F�w|�U�G|��@�R�>?�Q����&�UB #�|G<��H��B_֫�۷�5X>�0a �����!�˖�����VJ�P>Ko�9n�С���3�%��W֬�s"�Lҋ>�9�J�������&aI�f���t�V�"�n��D��3��n�����J	J)�5y����Q�M�:�1���D��8��ʑ���@sp�ѣGK�����4�;�B)��lU��2��=��	���	Y��f��Q��@Kcill�FaT���2�T����B�Æ[z�ȕ�6�6�by�Ȗ�P¨�
�p2,Pưj�8��8�1�;@�o6<]Fg
��iĔC-=����h<6lBm���WY�Q�w.��ssk��Y�vc=��
�#�V�g!�����}J !�	
1����P�����(-7��0�1Ɯ�qX[�,�%�N�t��R���,���Sa4�b����w����'(������N��ƌ�a�g��T]�*V���L&q�b%e*�c�̻����TN�3���cdRWHii�T
������N	�ֆë,�U>T�6<���ca�ň��>�MX��k@&�8`8��555��Uk;�1A��4)T�P�)�k��4�݀j�ݰY	4Hdeeɤ�
b����ʔ��2R=+��r)Z���f����x1۶m2�he��ׯ_��X��}���LPj/
6��P�f���~
�8W_�c@�WH��̒/����7o�,C
!�IOO����	ci��n+��P���UکS����Ƣ���ۅ�����Ł���0	�6m���K<ً$�ݵk��R���JVc�Q�ԯ[���
��v��������G����ھ��bYYY�5��]�����͛��!�?"@�2c]�$�PE��D�P�
�En�ym��N�/z�������35��T��������s���S4�l���f��r�Y��W̓^&��B(ߏB�`����G?�%��_����Ez)|��M�J�4��D��.����ŧ.�B8�6//�h��4�ҡ���R��C��q�j��J����5�G��ّ�s654o��ish��J�YW�^m3f�^�c:�����"L:}�Y�_���9O��z4d�2�O����O ��'\3��x���x�-�?��0߁Q�f��$��� �JJJ�V?
���wϕ+WDo�U�Y��B�;�xIxK��@αB���ǿZ���+^?O�;yF�'��\��u��?���Sxh���)	t]ߛ�_�'�S��E4    IEND�B`�PK   '6X�� �f  y�  /   images/96fabd4d-0b16-452b-94e2-688cfcbce531.png�	TSW�6~q�i�2*VA �Z*((�'A�0I�PQڊ"��"2�A@D �A���9�s����������f-���s��g�g?���^��ݕ˄�A����F�<�-Y�X�����_>~K��/u��A�����������t;�d��y�����)k�h�>s������mĀ�0m�j�;��k�w27���$[&f���tt��,�ｦ���ݒ�_n�1�`�=��k-]|�!so�O�~oy����B?I��l���K=�w4��؉#�[^����c�}}҂#n%�@�'�M}S�L�d;vg�|\������zƺ�WOڪ��g����VW	@*<�6++KK.��6��{��4紧���;�쇿V=漘5��L������9/U�c��r��;]�[�Ťk)�zj�]i�19I��DU �ƻ�{
!�w(;\Q4�_v��ͪ6��![�V���1���|�;����0�j�t߮9=X0�B.���L�0�C
�17��p�d��ۉ�� �n�=]>�����A�oVtɻ����1�Nj���v�.&F�3T�gČ�iL��S\\|����7=5��SK�����,�2���؟=���/ʖ��k�޻c�ׯX�p�@|TozƬ�N�Q�TcIx��z��j��xd5���:ﭛ�_��cz����5��V���D�Va	-$���E!����Z�����n�\6�^{�-��0~��ߺ*y�MJ��_����s�r���0�Y&Q�wNउLL��V8���@�%]�A�?���z"᫇�\|G�*�ς]��q�����"�"&"/��M>&n{T�=���j;��{#�-���~~~�ѕ��Fd�UD_��a7�rQ�2�ۇ��.M�H��-��y29�H�Wwg!�
��YW� �ѕ�=�QV$_?�l�m��7s���H/ds{W�z���]��Z�w H'z�S%\���4����_$����Lz켣���y����a����vD��WU���u���#0�O�qb�П9���!�������@!����^�}�{�1�sN<rĂbH���Y\n_��e}�NM�*l�1׀w95�����k�;ga�<T#�B_��zu��X���|MPb�[{��O�%ot������$�u�B������)ڛ:�F.P�9����3�4���s���,�D��Y�!I����I���0\��4�����2ښF0�K=83�jLӐ�OV{�;T&���{6��mr���n�9��2�fq'.�ZҜ=�l䣪��5��9/���ԙ�6���y*�w��,+%UF�lr�M2�]y��]4Y�)ˬ�ޅJά�)N9]��� SD�,���.����^��<7��]����))t7����|���e���\I⤌�p�+�4�m�!cE�Tc�ۧ��O�����`���4��BO\9
����NHk��<.Cȝ�#i*�y�YMMMK�,9H�l~}.]�c�����86VY�Q�榆�,���\�Ǉ:$bBU�Y��A�C*�dz�gHp�x��)q�8�;[� 󰱝��l�W����\l�G�.��+wI�l}��v�;��a
�Ӎ�Y�wVA�x�˾�h��&���@{@����ւ񕒜9KF
�-�:�U��]�V�ç�2�ko�sn��z�ah��d)����
��mN��e'*�[�rFXOX6�[�D�ħ�!L�iG����I�P�qT�G�}}���{o0�N��s�x"����Y�f���]�<�RdX��~��cz�Q�t9�H-tRv�H�N��=cn�a�f��fk���[��?��B�eΉ N�]{��&D������!]��Z�=q��o��e�~�8'Os�{'������r2�p;�CD�zݽ'i������܁�---�=���>�|� �"��5�͎�7B�=[��_�K��΋7�d������f=N��s�����0-]K�S\sXˁP\uz�����UЉ���4Y���xM=�yp�A�s	-b��wn�ϻ^n�34W�pc��Y2rEA�.��`�{C^���;UaG6hsl��)h�(�Є��G7U���d]266樫m��ކ������=6z������-�Xw�a�z�Rt7� �$�](�B���-��s�G8��YhU�� p��r��v!(e21���R0��~��z��F���VnYM����љ9�tM6{�9��iͿ��*�&#A�o�g}�Ɲ�q#6VL�┘ds_��$J`����y:o `��/wti1c��?r��m'^$m #����K Q;����ֱ{��1;J�uC0�0�{��v��h'a��a̧QJSp��W���=���{ ������q��"-�l6ȗ�2  H��f9V���
�K�ȋ@�h�
 �d�W.��5r3�{k�Ó�p'u_�"\��F�V��F�nz���CF�����}zvNMu��x4��<�5b����Ҩ�,ض,���R��˗/�2^��o�a)�\�X烠,��O�\	�����*�W��KJ���a'��d����H�4�%�U�Y_��DgK�TlB�m��E���iÅ]�Hٶ�h]�� �T/^$R� �d����X��\����^9ɪu�uM9�![%� a���M0fJ�3�:a�f��A�8,d��h&���X���dե�fҔ#ybvz V)��R!;����2G��[�'0B#Y4͛s��ϺC��@��l����N�.���� A�b��(��g�H����\U�r��ٺhONl�Y����K:�
��g��ӱ��X��G�Qn�Q���Vu�ƾ��0�CzL$�%�j�M��tG:��|�2g��_�����~z����' ���p�R��X%V7D|f��fx@^�
Ev�9�jN1���v�Td紊(pO�#���sl�T��c5��B���Uy(��&�)S��&�\�$Mw�s�zn>�	ZjêkG)��=]��wX��JQǖ��������nE�?@j�����}sa�
?ᘗ�i"H��	T7o��+�6����(g�׶s%[����圀����DS��Z��\���y(Nz�DO1hXaD�J8�\�����;w��������,É��6W�i�����e���|�>�@�	��6��M���WC9ɵ�o�3L�@a,,͠D}*I}��4c�r7Ǖ��cNZAn�Ct�ׯ��}��u��9i��
�R�B���qW����Y|��i�κ"��ۦ �]p�o��	HJ�;=ҳ��8��1�*Q�t������p��q�^9ȕ�6]����Ɯֺ�'�1tqV���"(}��H��l�0��h�0�5.�RO�_#�#��gPrgpH�f�z��`��زT�c�T��$1.��Y�( �(�t+AzvI���)?�hD|I��Q( �
++��9G��G�g[F+~����&�К��f��1���g0���G�D�t�jDG�����E0��p�S�}�]��-oQ��=BPbӥ$]�n����E�x�E�.�R?�Y�CN��k��l	
X�É" �XM6�����q&;�Z�`�������D�~w	4��<q���J�����uϩ2!���E�5��(�8vu_�q�qL��5���V-; �+
��cb��03�E��w@ˇ���1�̠�&5og�;8��9��=�N�Q��(�q������H��9 �)��|����ŵ�#r��Ǉ�z���s;�EͿ��-�PN[���Q�۶�:xF9Ҁ�
��D�x<ݲlf�9�W ��xމ��=)�<ǀU�_p"��0T8foZ����Ć8�' �U����3�ј]s" /|ŵ���6��i��F�Y�h�֊���n7a9������l����52�X����zw�0�T� ��ӳ���K`���/9����
�N����
/ւ]q~�4�ڠ���I��R�zU�R�%>�`K�e��@%UI����_������FI#��o[�z#9oҽ��w4h5�o,$�K��úW3=^0��b��'��պ9��՛���'��A��[8�����֒P���\��
q:*��WO�����5�Hl+К���<u��l@vyV��B�(��A)�ưi6���WC�����6)^�� <�]�T��:�E�y�K��DϬ�ǽ��5��;��_�ѳ��)�N�Ɗ�`�p�Ig�(y�n ����|+v�S��J U��)�q���g�H��} `��\n��;�C�<�����Xxt���,1��;eJ,��-����ӢI���^�%ڍ�j�oŵ0�mn�$�ܩ��(����wS��QʨfĘ%uf�t�a�ujR2�H�tz�W9*3XSQZ9�7A��W�1!�?#����Z=� T��'_���vd6��`����Y1��y'��;�'C����r�[΂̉FrD�:�(дTm�ZUcBgᓽtV��%�Ŗ���m�����55����mQ2�����sYuM���~B+�u?���=��}"xl�7i�#������I<=��.)�{�z'�[Us@��a�q�Ғ��Y[Q����I3Rr��D�O�ƺ�61�LZ�<|E�Z�C���2������<F�`���F��֚��N5خ&�^�w�	U���:��٠�Żkw�ZE�\�ʐ��w�����)}�	�j)��Vs�ۊ��X�ЗFRfӱ�3-���{�zb���Zw��=���͠���(:�w��v��qqX�M��|���-;������K��֖K��I��YV� Zi�q����c�|0q�l������Uº����4@�5D8�i�����6纜�B����pŮ�D�שr����錩�<�B�Qf1t���Hm�޴j�e� XUL�b�'\X}��O�
L����i��olA��(�2�~$Bc)�-�9#P�����{3��r�t��mS�#������Ps���D�΂��h6���ޓ��y��Zzv/�(��^Lb�^����0؝F�Q5�3�r�ӏY�)��S_���ꝰ�m�sCcb>`:^�Lc�b�7:ekK���=Un#/�
�zk<\Yv(F����X!�{J�����zW ��t�s����\ˎPF�/�&�(�&Oh�w��a�<��6��B�1/�'��ş	�~�rl]���0�����oA/i8��lz�E%na^T���dd
Ut^q(���M�����-�̸Q:bA	z�[C���;D��89�0�zq�!�4g��gf|uw�4�4$��.�I 4�?;[�Y��[8���9S�'�BHjH����b�pؚ�����T��1.�`5f���KI�YWԹ}�2{�~b#A�h����2�\<� �20�VۖA"v�?7�ۃ4�"��������iP�p�"@�a$;�����}�*n��� ���d��-��'���|�漾����u��ɬVKJ*�I"ܾ�Jr= �v!n�r�!�Zܸ�Q���D��3+'KnII�����(Зc'��1�"����e�
�o��0�p������d�.�)� m͟��H��#�K�9�%��zO�nS���Ld=2�1�?���<k� \�������y�����%����p��� �U��[%��g�V,�¢��m�Ŏ�Vg�E�:f�W�<ȭ,"Qs����ÑFk�څRh����9h\�*3����������p��t��|�ۛNZ�.S~;+��p���bkc*��|F!�=*O�M��nM_�B�����󲹎���[W���tC�t5@���d ��P0������
*<�L�;U��M5���q`}�/C�p[�ji��kd؛yy�C���`��$�S�[25����	��c�Q>�h���\��	�t�	j�{�Y�5]�<�y����5����� l.P���,�䠔�f������+�\8-�p�-�e?A�b��d�"�(ǫ��{u��#�J6]���pݵ�}Z�� չ.��8<�b[�,�&�K�`G�+i�ۍU۱��&�'�-lϗr8iP>�A���P軜"��Cl�-�ध))��+�A�͢�;����,��tfm!��Ť.@ڲA���y��w	p?|&��PG�&���ښ��)5�Pɴ0��&��r��}λ e6)5f ѪYط�� �0Z����p{}��v��!���[гVШ�y!�;hY���lȲ1���y���������"e~����Bз�M��:K��������էxJ�3�Y��G�WB�@��P�IF��L83�cq
�֜�.*&����0�lH��Y/l� m!hi~mry�nZ�����iƞ�2s�{�[8#]����&��2{C��y
j���h9
�I��!�f�6�O��	�=��(T��^7Y�X��i�sQ		�:��AW�ú��d��t�v�%姶9�B��ŗ�}����4�~��s�) �K�,B�_�U�?������qnv�m`��ڠ⎱c:�+�u�&���&^k�MP�z S1�w��jȇT'�A��m���|vw�jD7�@O'n��o�VE&�8Fy�+k>{�84�Z��~����������?9�l���;��^�����џ�X��	?�M�!Yǿi�㭗�s���2���Xq�R���Z�^u� �hB�}z~)��14~��F(b3�\�e�M��W�p~z-`|�&��َ%�X8W�a���9�'@�?m��9���Ț��{H�A �-���7�PkVw+ڤ�O���oHӒe=��v�%�5|F�CŬ�ڒ���-Z�l���=�A,���ه`��S�X��<�ۛm:���G��}�ټ��=]8� ��N�e`IU�l.��c�hp�{����e�d�Ѽ�A)p��[rΕ_X��W!�����W���V�
o�ɖW'r�n�r22�Z_�o����<ӣ�ـ㇭�(ہ�ey��.�>aN�J����3S36t������cT�8�d��j����$P/1�P�Sߩ�4-v�'sȮ�CB�PMj?(�0'�����*e�R�a�l�O��=�l=���I���
FYb�)K�sO��t��؜�/?���d��G�il��ϒ���䲟Ӓ9�2u����,�E��s���6\ÏR�9���}S�{/��w	(���cЎbG,��/猋��s9�+9��W�c|�{�B�D�N)��>@���:9�T���s���J�ka= G�P,(�8�����^��~�I��f��ps{��w�����RR���0&y77�n��亨D�iE��7�C�i���&��@u �:%I�� 2>ݸ-=-w>���I�0ψ$�^����LX��x�3��M��(I���@+�J�>����Է
�Y�}��wKj�9���z�Ϧ��x�շ�2�Bt���
}�����ث+
j6�6��!�#�c7��ى�YΏ=��څM��*�s�������[R��쎇�:�Ŏ8'���|O�w��ʋ?���z�H�<9�:r�1*��ͫ�Z���K��&�{���~���bK���Ǣ���o���t��}��I���~���r1��M��BC� ]����z�s���4�� ��z蜝��J�L�}H�5I\p�N]e�U4CZ�f1��cvGv�4��c��B]�i���p�->o.��fWT7Թ]�vmfˏp��.�����I��qHPCj����HS�'�zqv�.ǷAj�}aF���J��DχzAW���n��j��9���d/����;3�j�H����<QA@��m^�΍�M�H3`�}��I��̦��ר@�J���ũ'XW��Y{��f�|`�=ˠ��t���-�2�r�`�0���F0ڌTz�Qs&�9����T*���A�i���=�$��P�ej�������|dl��qkAzzd�>�tU�4(Mk�48I�4o�Y��y/�GWg�]�Vp�I���P�c��%_��Ž���&���$��N:�ň��T�f��x0.�b�َ�m�Bo?||�l��Lv�fsj���q&j�2gaFeNP.�3-=E�PSS[Lu��el�x�U�G��}������e �؃�<w�r{g�-�op�q�����p��н�|R�*k��܉�Re}�n~�.](�b���"�7��΋���?��.�A�n�ºu��Gkf��0�ys$�ʻqL�UEa:��^_,(b���`D�ǰ�@^�M��\6�V4�xyqJ�!��Wp�R9i#����%��Ka���?�q�{��� ��魷�4�[����LQr5rb!�gÀ�n��n7���RDӅ=�,*㤪Ho3�7wgL�|.�(�0���!7U��`@|�e/[@'bz3/��2�Ҧ��ϑ��Nn��������j�R�c��p��>q��#c�hE�=��_�@�Ϊ�Jbe�?YPn�R���K��Ka�$W���­�I@90=pYP�+z���ƹ$Q�����J̪�Y�Kf��Fֲ^�dj[J�fC�K�+-�����:r�=P�r����Ĭ�E�=A[�eZ�P����]��4�pJWH���4LS9�49���5)5W>E#~W�A�M��ܡN�׻7UMM&�>�P-��X�0�q*��~��k�'��)��^Ajj~�D����TMu)Y04��4�`�aq����Lſ�D���R*���rnQ��	z&P,�=�������{�#���H�$b�@���&gS������1S-gf�Dʞ�	���]����	�������=�d���\�?�n�����������������������������}�.&F�?i��]��@��=�ֽ�Q���u�e�˙а�K�S�={����L�ym<�8�+!��B�qO:�;)����C�#�7j4G�$�I}f�M�K���`eb�Z,�G����#G2���F�&��뭣�X���!q�挽�~(��F˭�	�k�*�����Oss����N��9�6�����V�xa痼�����h%��Ω�FM�P���ƐK�ǐ����hh��Y�Sk��Sr{�ݛ{wwe~�c܏�n��d|P�b�Ӓv��2g�<��}�NIL���=PlK:�tAe�@��"
�>�u��3,�,�9)�QnsN)"rʧ������gML���ه�:��z��?��r�������q�/�i΁�w������[��ឍ�>���q��7�{�_ޘǬϊnR	PX��P�;��ҕ�5��+*�eC�N��]��Uי�{Ϸ�^�s6�]��M��-R&�:�7��5%;�F��q�2�e����%>����}��,�#Ci�}���K�����K��@C�i-�)�c�=�T�;��DȐ�9�aR���G�a��C!�M�N��f]�+�\�Dy�vf�BH��$�B���ֶ?�2�);]Nz�KIj��A�N�ZagF�r�B�i>4��?zo��Ջɋ��v'�F������
�Yu�+�ϔ۴�T�MLu��qvf���ʨؤ���x�>�Ŭ��
���{&�Ns�������� yG�@�|\\�����sg	��mf�ŏ��Ë����@Hq�G(��άoqs�e���h2G1����K��GK�Zf:�h�9��b�r_�ϫ����l�a1��!�8�}gggBL��p]�&��o����dd��O��o!�����	����@>6��M9�l+�R�r���t�����5�gI�Jc��������[S�\���X�i��
�M���*؜����
ͬ����
��DV�2��Z���di�(Qa��|��+�_�ϑ���b����:���w�����
c]����'��`��8-D+1���D�l�Gu���t������Kjy�ZӃ�}G{jz�C��`{Q`��%��x�.o�l� DX�r���	�%kwӠ����?���͇�z(��N�2�A���j��~�]�r�o��SU(/�'̤�ncA��:�O�Մ��?�*[_����G�we������o�v�X'�
�p�W�d��[\ބ
�( m���:��g�c
y�Ajq���%��M<��'�D����@PzJsV�:�^M5َ󯣃U	"ZZ��*h#��"���V����+)Dg�!��h3�	|˸����0V�2����*~����KJ
���R�k�7݅w/&��W���!������);!����
�z�_�m6�H�Z_+��n���λ>"c�|�.T��~.�kV�
���Sn�ŤƗ1�m+�Gsn/_d-7�R~9�O���m6����� B[�W]��-P�a�"�ٯ�η�a9y�u��-��6�\
Av���< ڴ�)WZ[F�y��4�T�o��b�_���	��#���ԻF��I���_�M�v3�k+ hծ�ry�ҽ[ѓ������n"Q5����ȷ���`�5�Q5���*��� [1�?j߻�Y��'���%���m!�91)	9����k+�P�"\�[!�{Q�������󡽚��MX�5��4��y2�G�������شC4E%��'�W��dM��J�Mc����׈ VΡP�W� �y�J�G�,fm���W��M����u������9���+���NP~�
A�G�w�$B$���)�������\�OW,�p~�8_⓯��_������_S�(T*�� (�%o!W� #.�R���s���t� �����s�x_����A�'`!���L�U0f]��`���J����H+㚗��w���S��.�<m��$�L@��J�t���L�"3��Oa����(*�Ȋ�����&����Z~��p	Xi��1 ��o�C�_q&���tij"h*[P}��FezO����X��r�K�׾_|�ja]���ѻq�YOц���.�:�A2N%�hVs��}�]����C��T:�˯*��O�7\�3E �(�ׯ����c�������t@�D<�^J'�9�Ci �<���V�G���ݹ7��U��X�������j@y���`<�!\��^� �C��'�'L���,�OM޺f�B~Ś��?~h�s�\{��|1��,�������pqۨ�H��0N�/@�t��H
=v��������d�"���[�������߉�K�|ʎ�?��Ż�F �EF��o��q��0���x�����5H�2�}n��Qa{/��R2�Ex3�>�+76�{��͡FC��ٜ�����2�U�?�/�����Ĭ��aS	��mF�N@�vgtEL���7��B��������� �]����߽�;����Y_��qtnػ���@�j6,�&�cU�ߋ�'^�k7�s�u_OO?�s�����Z�C!Z�Q(/n?���ۡF�w�&�nE͗M��F �J�Hg�{��G�@{� �ٺ�3��2�c�V����$�T���~c��@���>�6%%�0^W�r��k����ZS��8�oK"��NI0�`�ay�g��Ъ��o�}�n�\�6~Ϸ�M�!����Um΋i�3�+K�c���ʓ���������T��K
�廇\Y�;�����3��-��X��쒁��ݠ��������� K��ļF��l�H[�vgj���;-�(�Z��˩��wF��b�O��t�(\�14~9�z0񋔆�`���hW#�LQD�y�����N��
���o��maN�,5������6�@Z��ֶ������F>r�?;v�I�՚��|�#̛�M��J�
yvƆ� Z����L�]�l��i� �{��z�v�����V�N�U`@j�������s�d���J`���L�[Q�\��Z����3�B���嵴�g_\Ӻ��������hÞ�وЪ�H��+Y�<ˣ����$A��{�ױ��ة4l ���Q~��I0)z��#˿V��n!�����d̚���4�G�k�>��Ą�ؼCQ<8ǅ�����k��	�P�v�p���FLL<mwww���
�L!VXQF��-���1���L�]�r�H��5�3-h����0�.�5Qr��~D��Ԯ���դ��2<~8'9�����d���qu�� f�y��WA"fH*����w�&��.����s��!���ҒJh���ҝ/Ȼ���nnktuu�g^�#��_/**:ii�y�E$�Uxb�S�V�M����
�� edd0��>uq^���`�S���0�1!1������G�L�ə=[5��笉�/�_�bl+�<�=ݥa��h�F쐕��W9�p`pql��
㔞]݅T��6A���cD�HL�e��f@Qnb/�콙���i�)�!�(+RE%����^���%��4Co��j�cZ�OƓ �͒ͯY6W5�V�vy�G�?�Lu"�֎�y*��-4ճ�32���W����H����Ļ��&�����Ӵ4���w�?o�`PA��;:ć9(�#{wz?f��h~���
#�j�/��a������mll��!�~��.c��[RɕA�Lv��v_]���jޔ�������y�ӓ�!#<<���f�u�N��ț&Ԛ�e�g�P����X�)��4�_�!a�F���>�J`NS]���79*'Zd�	����Y���b4Pv>����������Π��(88�د]Y����v�l���.��LF~�g�_�g"��]L\�Um�	��������L��7=�Z[]]���zݲl/ě"I�I:4����W�^��[=��X���'E�b��3�+ ��V�T�j�_���N?)���c}���p��H)"��x�ԩ��1�'���J����Qߏ�۠P��
��l��ɧ����Jt�2rժU�Zr%V��°�����'m e�>�s���:�C�{��wQ���]N��	i��W�H�x_JE{J�f v����������>��Y�)fć<a��(�3�n� i��6�b0���-*_Z�����L��kaD��lR6DP?<B��mI��5C���xQ#=���. RGc07I#���*��̞���-�Q���>��(
u�А���^&&5����3^���Ky4@����D���c��@���=k�/_�4=��[v�����Q���Rw�Naˁ�,Đ�^wf����&S�<�.^L&���i�ɼ�� 0�$Z_e��]���]tfp��;�HT���5�t�>�[���Ei��#��.���(/+��~� �w>�Ԗ��Hۜ9�@R�]:^� {�d	X��4�1И�B�5��I'�������X{G��\��Gܲ��+
[e)})J�|~t�p�ATDdd�|�,m1L̕�N�j����d�j9,C
3��[�̙b�SB����]/^�8mo��^��99]�(�F92�%8 ��T���]�� ����ʾ��m�+<��`�U���3S�/F7 ���?`hU ��ddWWW(S��C�2�6e���dV���T ���Yb(TQ�=�Au7����툧�e�ff��U�ώD7�{�	����j�5xO����pU���(��熝�K h�v>�lc3u��G��`2ГYY�1�K�SBR�P���xt_Qs����P���� 1�Ԏi�=B+����x'���
��#�1�]u9��b�mB�s�$m���@m��'OΧ5Tv����NH茏�$�s��Q<}�Jk Fh����L�u�2��1\MD?'���m>$�2P��<sr'yy��϶Q��4�@S` �*�"�s���'��3�)�M���Qvt���r3��K�ݵ~�I���m�,��cH���㴭����{�D"�B5�l��)2qqq���7 ��D�@|R�V�]�l>;ҥ��W�*4B������J�B��R�v1I �j�ʌ0����H��%˭ꦬ&GE�$�#����c0+�<��%+}�w}��{|e���T#�Eu���������⎺����I	X�?
�	�����5]�'��0��y889��O�i*( ��Ў�	�5�kIꝌ�+C:�Lʹ�z�e�ڟ��@@� �XP\��)�A���T���Mh��l�� e P<����#0�?m)�(,Wn��0s"��̍<���l9�BT���p;��A�&SR�y�f2����������u���!��S�"�\"Q<3��,���A'��:б�o����M�(7ZМ�6�цdp�L@��Nar�9���BR�I$��xG��1��,��i�^7 vy@:R8h�7s �:Wr����cE��y�e�>q�y��S.��5�;/+ �OĹ���j���a�n;�]�����qfgh�v�� @�%d�Aѹ	���$��E�]<I�����'oe&2�^�d�=I��T��x�g���Hs�pQ�该21��xV�i6f�E�����ˍD��"a=���Ǡ-�*uo��BG�,1�_PP���~󚠄N���!"B�Fjr��N�|���Pt0p7�u+�$E^Aa5`)�]P;�aeb�RS���u^�}Ro&�i���EBi����s�+8X��+B�l9��:�:�'OI$����J%8SZ&	E5۹�?ाLBL(�e��i8��#c� 0|�4�[��� ��
����n[�-�ߣ�0�@��Q���R�*�ng2�i ��=�|�_ ����1A_Q�O�'�,-M0\�������ݻA�Y����M��D����쎕���&��清���/��F+���L��N�N�Nk�,--����G}í��O�4�=P��~�W����b����ک��z������9�&}}�����ޢ��;���;F��23�{�XR�fW�ׄf$xN�:��ȶ�ZO�	�#\��5�5�Zx�$�F��Z�Ύ&E�\8��/�ٔD ��ڀP֍��XP�����^��B�-�>u����A:��ҁe��I����EnG�b7���HH����h���G���roNLL|���r�`������_��i�SQ��K��u�{�,�<�LN��&��&��=�O�@��>^��3~Ƞ����quD�z���ji���O�y~�hr���;��&Xao�篵��C:*�u�}��$a��<���/_���y!�6QX����ud�&m��REEE���M����?7M }w0O8��,���mx�>d��a��W��;
��O����jۣ�XC������8��sF�u���Z\'��E�4қm�9IF�Տ�@3I�o�G�����#-3^y�GQew�p,?�$)�\�?�R��f.��F��J�:L� �_d�7\�ag��|��u�C��l �<�a��k���ƺ������5�6�ު�ݱ'J�.���U���?�AxC� t��m?mrǋ�u����(˓�^gl5UIA�mf���	�?b�)��`g&{��t,����1*�
ᎎ�! 2��I�Ɩ��&�l�̤�V�v�!b��l1�+K�2�<����6�0ةP�8��l>6��>4$/.!��h���r���9�"ch��a>L�`X�񾊢t�gq���4�l�ι��Nͅ�	�YK��h�V,oHC�pe1�v�C�ձ�m��A�w�����o�\��ݛ%<Q���5Ђ��/��-E�K�x����CԧMJ� ݵ�ӫ5w�W��,:��>o]xw_��"���މY�V�s�BS6�$oe�w����{=�'�n^z���\`��T��O������K\a>$���K����S�6�*�yVI�w�����z;�	��[���I��_�w�o��_�^���;+.��m��χ��R{��@�%��!���=<��7�@�%��&�D�'�Hֶ�6�F�M^��u����:��c��&�/?�ٶ�f�N��p(؆����<�p��M?��]]j��}Pr��dYQ�|]�L��3|9r9��>p�0�A��7X�]���o�y���V�q�+%��ٽPr,��!m��v-�;�+[y��~��}}�K�1���hyz��H�8^[#dd������@�ٻS��9�`��;��Xx��K�hn#��_�� �;��ut����g@���ŗ/�o����n���o������?yA�)�
`%<�j5kk^�١9㣹�-�ʧ�o�����@�������y��e:_�(S���H�O6>�9���Q�{�o
�l|Qt�n`�����0����7��pk��n߫5
��}�a���l J�������,d�8H�����AQ�V6Bz�������p�͍�]B
��y�������̳�� �̹G��_��S���>�_� �D�η����T����I\�u��
�S<^9���|�`:ߏ���D<�}{��.��W�����t���n�Z��l����*`xy���!6�_�:����.GȼxiΦX�6P�&D��� �� �V>쇜ݬ�y���0ʻ�kUa�p� �R��v�ڐ׺�K���E�������${������zo��m�|N^����9�	�9%�����d����ޡ8b�f(�[��{>�<���90������r��i%������_�q"��}1Du���'�]yf�[�K ��;ͣ���8�2�]f����jcF�c>���������m���"����W�8�Ւy�ڈ8�=�5� ��Ȃ�)J���_L��y�N�l�S�۵�l�w��+��ϠA��Cbu�^&@�':���qq>�G��?jȤ�W,){]6�4��Y� *��V��&N����J�q��:=��?���'�x[DӏM�z��������Sޔ�{H]}j��"��_�DxG�O��7W}���I�Mkxt��Z���ew7�a��eu�M�dRݟ[k���H�o��}V>e֡��#��>6�>���ҩ�oӾ�<=�b�J$�M�K�\�Z���?�-z�]a��I�(�y37��{ץT�d�����W�/y3�
s%N�4b����t��<t�|�v]
�����F���TxA*������'X�=x�ܛ,�k�ª�yi+��$����a�û@1_AVm�~ H`�O��N�C]����G@���+@��%ށ�>AX���ޯ��OQ 9�Lɲr0�ｚM�_j\>S�k��9�|�h�I�d�����C.Z��2����]�{���E;��}�e\��L��x�!�BGy�h��s�T�'/7C*�G��Nyx��ٞ5 !�/��|Z�Ma�B����ޏ|�anT�2k��	`��_kƹOk6���n��G�V�/��7��b�~Ee�E����BC�WD�����^�ֲ�����6��{���5�������ξ��(��ln��	�D�1�)t�Kl;i�� �n���#`�Y�dz��?g�����
�
c�ྔ�/�0��/;�?�$��l	۟������ѱ��F��:�WF��6O='�k
l7��>�d h�ꗐڕ}��_l��f�����>���F�<�����u���S)�ˤ�ӝ��!��Dj
PsC醹��x��E���A�;�8�v�%�JA�d��R��
�9zy��ҳ�]���s6�������r�B�~�<�q�~����O�QV��7��9��&@���%g*����kW��]���4.��a�`N|�;�H����~��$���?�R��ħܠ��k���̗��ؿ�� �`!�,���aF.�ka@�#������O�#> f��Z�|E)�t0�%��o��k5�8��y|(�{�<��I@�w
�-X�wun�������X�c3�e�[�~��蚮��� �u�����`�ξI�d6�?)楝����@kp�Rz��Z9��a���p�n=���u�m�I�<��|J�<�fėg_��{��F���&h�=�hp�L�.�6i1�d�%$�X��_8���k^,��ټ��4wp��#�D�R�~#ZkK_Sӯ�T�!jx�@��x���N�n�j���7���OF%Y��ɛ}�����n��Y�I�z��/;tm~����ͳ��̻��:=�҅�j�oI�� J�L;$7Bc�$�"9� ����ePF���������/�i/K��x��}��ॷ��yn�,t�H�BEb��%^d�m+Ux�6�$��>Il�>㳑�`d�ʁ���Ep˩���v������`Lm�Mf�P��p�|_�/ ���\ܓ��a��jcjƼ�!tK:�,vh^Ŷ�f��E��렬-<�yp⣐m��˙�C�3ߟ��yK��лe��������c��릿Y�=@)�;����E��N��'��^��h�)�g�~#�Ʉ�yG����u�0�^i�؃���ޟ��y�zA�YS�����S!�ao�M��"g�`���P��= ��2?��o�f�f'[�m_!/a�T!>�@�Ύ�y���d�O!���yq��Tw;�W�Z�my���������%�E�ƍ��;V���^�I[^_�{��7�"�4?��K���͇5��W1.]�[�x����0�##F� <{������i[>�v2��G�8�jp%����+��L����?� ��\�>���W%owT�j���/���[x@��h��(�X��J���|^�_�P��%g���(���3��?����"��`^��~��:�� x��ڌ�}�}��ʁ�+x���A����ὭÈD��b�4�[�<��e_l��ح��^u�oc�a,�3�u�N����	�$~�XO����!/ю!��
��x_,P��.����Vrb]+&u��)�Iv�/�\���E����rd�A�L����ѕo�w}�3=Q�44���dU��F�
�8/b-��$�<��p��[�����d�=������9��^�� �n�)�R��(�Aޤ)A.o�8`v��|q�fq��{[�D���$F������Xc��O���e��߁�F-(�G}-(��	�-���hM�{]�����Q���F��4@G)�2��*?�(,��ur��Ҁq��h^�&����+~wk48uރB��{�|x5
�0�6D�݀<�Z���){�oY��DW4����6p�{z�^�y"������*EVkw��/Qhƥ9\H���xx5ۅz�.���3L��r�ǝ���1
��n	����:�n�Z])��������<��X��Xq���!͉I/����R]�mGA۠�1�j�^�	#=e��Ս���>�I��8e鰵�b����L�2���<����R��dHJ�.�^�Kʐ�/D�e��8V��x�8�j<��{q�����<�/�E��T��I}�A?���YE}���G&�ߴ".�DW1��4+�dm�>��+��ÚJ�}csm�ሂ2�� ����r���$�"�� (�
���Ƞ�AeN2�`��9B�H		����>�{�}�{�����^��?ػ���Uk�֯*U��!�K�|�>���u�O|����^������Z��OE�8&-q�g����`�$/��UJj�L��I��X���/r��
�3�Cف�[ �6�m�F�.J�(P*�;�Y��h�R5�W�\">p"���-�0MEɜ"������K��݊����R�1����&��S[s�#w�GB��w�z��p�߶�ZYZ(y��q�q�8�eu��9Y`1�w����p2Q��`C#""���1����o�#>ǳ�D��Rֳ�9l���r;�*P9� q:4�i˥L������5%��@![�}9�&����Xÿ���}Lx����<Hv�)_N���6N�7�(��^ڑM�.ܵ��뉫dĤ��ޏ���q�<9���=��)��Q��&��K*�|#�i�S�c����%����_�R��9�k��M���Y���礪�+L�� D��7��+ֱx�s���%�������	�m	7Ʈ�~@^����D�$!����0��7%�3*"܌�����Y� .�a����~E�M��`^L�G7�� ���)ϛ&(��t��|{�1�#[�,�6��4e�����z*���lI�����V֚�=��V��
�Z���K@E�u	X@�oR�&[Q7�(�V���+u�P�5�<]�����J��=�Z}턆5d������9r6����b{t�AM_;�߿��i��V�Ujxyɸ�S������ֻ������w����>�I�AG�����;l���$��`�)0b�ʘ��ϗ�T�M��2T���@��W�p���D�]T'�'�T�}����M]V�|�*L�^oj��$�Q��=��7�U�1�r�=���!�����ʈ�2��[����I�'Na���-��Ũ���٤xg�z�����g��U�7o>��Rf��j�Eǃֶ�k�y�'E���`���/_'R$��f�A8(XhX�L��Vg[� ]��%/�Lꥬ̮�T��7x禍�i�/��b��~U}���0p�&'~����q�Ĥ$�TI����@�c �c���P�_*��3���B��*vtx��X�WK����b��a�j]z�������vk�u�2��yy�k�I[ 9ΧW0�`1G{=巽�o�K�.��Z-j��U��`*�`�*ʠ�ƛ�yܰ:i %����L���]:�%�ɐ��J?
S�E	��f����,�l��M�'��7e�Ol���>m���)l������N�eׯ�N��W�Lкk�ޜ�?}�����4��Ջ����tf��!5~Csssg�����2����@p��7o�H�D*�n����B����|�1��=�o5�I�M����%���QdT�ߺ�`$��볘��$)�> �׺�q�+K֋�L���*L�ș�Q���,�[a�p?zt�Mxa�J_���6�`��m:�P���"�A���Q���{�/��L�J~�?pa��5�s?�A-���G�'MB�`��(�r���`=�C�%�I��~�q}���I��58�����In���
��I�=��c�2�;66V;C:�箏~�FV	��E��*/\�/�h�(!����	��N���( ��R�^h8m�V�Zu5ֻ���?����=Xuwa��z}o���q����ʻ3�X	�FN6�N�q�n��(����3��*��'G))'??M��7ٞ�:b�J��������\�n�u��Q�Ԕ$K����+�-/�RR����sM�� t)m�`շ�r��įC;�S����K�%�g�'=�OYs*P�U�o�Ye�n�cw��s*	@kq������G
��V�I�A�k�wDM��%��0�B�ׄu۶��:���!�#:��J�_���>Nqʦ�I\�'>H^���#�7&���t{�>����c,���MMMSA����=����f��x�Q�%����P�Z��2B%��e����6#�l�hnz�p]:p�����s�-^'�%�g̸|e�v�R&�`�t����z�� 6 �o>�Z�����ܻ _I]�5�z~q	>�C"߮l(}F��v��{%�M>Y���= �W^�t~r )^%7�֑/	�}����m��b08{�=��>������Ѫ)�:8���*�D��Dݵ:	��'���_�I�|q�̊i��q�1��$Z���� %�D���5���lRMpP�	Z�_�	
{�}gǴD4�l1�=�3�(U`��OB����S�,e�4�T��	�jev�y�����O~|���(��c�5��.�S���#p2<�s1�[�!ǎ���D�� ��~�[�!sC?K���Џ1��Y����2�E1�PU�����`" -#�]?���a��G�ېW�� E���7�_����L�� )FE�m���V�޸�)��X�:EC,�߃-���ץA'���8�4F2*Q(˴|�?��#�M4�x��|Q&zௌ�P�N�Q��~����ba--n�ys'��*}	�|��ězg����vY	�(�@'�1���eC�����8/�j .�q9�������ݤ�AIh�(��(WG0杳�Z�A�g/����.�d	�$��1�.��ԡz��@�s2�`ʳ/*�5���V;fQ~�:Z�"��{����kP�� V�ea��a�ꞿ�̿����~����Q#ӡ��򺓐b)p`�`�P�fЂl8�ֱCPV9G(���hM�eX�[@T�G8ȫB/�A�Yd���}������o4fL���4&Y�f47x�ɑb���H��A|��(˳�f���{����luEb��(�b��*�ΏP��
��=CN,����+���b��RF�+ �d�I�i�r��q1�x�4gQog���{��S�l�'�;��8<,&.}��4P&�S�.w������I�X'��ʼt�-?
Y�ܯa�?���^.b�F`b�;qaf �o=
)�x�a	j�`��� ���5�����_�	�3���u�2��SR���L������/KY�����ԪP�\�P\D[�@�{���;?�׈l��������W �zc� �جm��2�kGA�g�wy~tkG�ڭ�G�[�Y���.q�r��zv�a�:��-�:J^����On��{��n��8u�Q�a�����L�����%��V5��ѡ��/v�Y^��"hSa�Y�#�x�e�g��D.K��/�����	��Ē(Ŭ��&�Θp�s�/JpM���Ж�^�ho���R�sGǑ'�!�A�����#�=J�����c�OR}e����+��ݹ��F#Z��%g�����wkoƄ7ekdtU��q�2�*����9qC���N�M��@0u����ʯs����JY���=�B}[w���??w$ԧ?�S�iA���y;�0�����bL}�>��+K�>󄹹��%��O��<0�Z��)��~�#���dۚ��V`��R{�����jT�za>��n���l�n�-��Ź��=t��[ny���|j!�?\g�v9u���ߤ�z��V�\h��%�ۻ�љ����i_)n���^��]˧��۝���l7 ��}"_��t��7�]����mK�8P��60'S �eೲ<و�#��(!��3��u]�Yn�l�v;��U�S�"q�N�[���NKd�(P:ҥ�����n�{�\���>B�����۟5�Bޤ�+��E!������'[����y�e�O͕�,M�;Yj�GFa�vlp�U\t�(S_0�r�.r�b/\_�\i5�ф�§ϫ�''a�~x�;�E�͠���龧gTc��t����с�n��B��2���oܫy&m���#���4����z�y�W�����s�����x�@���<x��R��y��CJ�	��s^�h,��P�%���sQ[���&��G�ܡL�*tV��ǫ���ݚ�:d`�~���ߒ��d�6l�Y��L%<��������v>^��������|�~�ͱ	xw_�����D�IYz0����X�=ٷgg+)�{M�P�)�qL��A{���Dn�*���=/�caFH��J��~Xٴ�����ħ#�"~ﮪƾ�%%j��[�@'`�^����D2^��d[c��@Ѽf�e��SS�������`�n)�:&�[͹������XI��҃���vS�^�g�� BH�����j]�Ε�N�N�c~t��^E�R(O]�^�΋��G���,7@�t7��1�"��}Q�j��z����5�Qx��$��Tp�K^ań��J0��_�'ʑ~�A�j�8N�F�z�d��e�G�y�ȧ����HǌS*OZ�;�W\������"�vnTۥ�f1������=�� ܋��c�V��S�(-�2Y1�%a�/Mt���jl�JĘ?�|���J
S�e\3y�Q�,�TQ��K���@jq�=�����]��&v䒾����鞯�������8v}��P�[U�ߣ(�=">k��f�߂Ѫ2�͝����N������ݮrB`�/1Һϝ`��w���	�(K��5���h!����β�X�D�5φ#�푫�r�3Γ����>S��"
�P����`�n�[XJ�d�ݍ�Q�+�	>�8NF9�|��H�qMۅBX�:?�D����%U�V����V�Ǖ��T���Ow.��x�\�����-o"��ӎ��Np�"��h�/�mz�a�+��Ƙy�f9	��o0WR����c0�	BwV�$�]���V�*��m�=��~���|s�j�/aV���+�h�͂�R�w���w"���,�|�Z*�c������\K����Fy��yZ@1����]6GU)ڨ�!-�#�Մ/"��������?�����ZU�ܞk�P�?�hmח%�TN���7��1J��/,,��'⸾�KK{�!�/�vZb�����5s�@�W� �������C������g��w}�ϝ?O���IY��J�����/�,?wH�ym����{B��#�[δ�d��kM3�gΕ+W��xw}~��d�G())��\5��֋pL���p*;��9��Ɯ�,�7�Y���&C�lt��p���s]�X/��H�rS.�a����%���$	���@uD��T|5����gn��OC�׎U�jp�Oݭ�΂;D"����%zy��6���z}'���"l0�n�^���|L��	��o���R�܉΂�߱E�-�}�l��3G$�;�w{�݀��c[��K��b���ӥr���p��Oa%u����'{RRR�	�$��mwf�B��<�P���Ca�����au
���Ȑ�A�ڋ�i|f�P�ѵ�Ę����|����H��T@��E�{��jk;̽��E�D/R��H�b�xOk�w�|81ϋZD�Aj�� ѣ=7\_O�L�=�'�)l<?�wTC\N�:r�1��7�`{��ɓ'�[�����E���f��3�-[���bC�k�����	&�(�|ľ�3��O�$IzQZJ�@�-��Oii���!D$��W�G�����a��偺:RC����OpZ	 7�ؠ��H�Ș�؊O�=�~���	��(���"�j
�=m��|���+�
�϶�M"��	߁�d��$	)f��������S�q���i\�~��-�`�r��y��ڍ����].L���r�(k{{�&X;�#��`��-u�0r�X0(�N��������e�P�(����lœuTu��oAh�R�����f]z�L���$� ZG���U#�kݽ��=>=�l�5�L���f��/���D566�h��ބ�g"Q���=����ݣ��ޚ�����EN���jp�77���J���`�+a�@�m�3�������G���Eq���d5k��UH�<H��s�v6��|�S�-s�w�ퟥ:Gͮq�дLX+ru<^�#m|��s�	��75&*��;��[�=�o�kD�����ve�$�]ײ f���9�6)�U�^��e��U����Il�>������t$]ۣ3�bb%�Z"k&�?�2�����g��X*A7�	'D9��

bY_���)Y���%�� Yx_A|!��;�� !GwSJ����������D�Ae�e��@
�:9C?�)�ޖ��������.]�e�p�,,,h���َ�@��Q�h[*p>7����-�b{�g���Ucŉ�/kdtv��1���a(*��PfFZu�R}���A�d闓����U���!�=ؙ��E���v��3��a��q�0#�Y����?�$	v���g7h�ٓ�D�5|>_` ��d1&'��}m����H$R���Ç �|��
''';�-�7��F�^��K�Iutuu�2��L]`l�O����eH���G���ˋVy�zb����W���k
��O���Tuh�k��i����]y1r��g�s�E�JIH���)��?�jS5�Z%��M�g�52$��;�o�E*4�����Rw�rLLL� 4Wfz;::bhA�,�1Mob^��[����?�ژ�pSo	*zC(�Z�kq����@=Ka�ь4=�2�R�ޗۊ�o��	
rd��ױx
�z�9⼟*R+�Zx)q���o���}���I���PK   '6X���5�  1�  /   images/a437e5bb-8d3f-4b3f-8093-72e2f97ca498.png��y<�}�>>*�,ݕl��d�=J�d	����-u�&�u�'{�ul�b,Y�!�1d��q?�������w����k��y�q�u]�����B���H���@�<�рW~;>��x=T�=��s����ϻ�zA _(?T��:�E���:n��~�6???!W'/+w!7O��9V�D��]���闉l��C㞲_��$⚟�	��eոI�OΆ{��w��y�V�Y��id&4K��ze�K�Ky�}�.ޣ�C k%��p7Y���:���x���T��"6��.��,��T^AXW��+���\��!y�Ϧ�U�
&S����6�h#}��c(����T�
Wsx��h6�c�B2W���k�w�Ht��_�Yx�Rǘ)��=������y�Y�	�!�k�\�?d��VS��(w���ؗ7g�usO��*��Y��Rc�О�\+�*Le����=>S�vײ����S!O9W1����@�k�EVS�J�Z���*��Ŗ�s�]��W ��ԻW�K�)�)�]�h��T=xϥu��}��j!�*'.�]�p�d���ic��:�k�|��E���c�#v�m��.����4g��~��t�I��D*��b�ѧ���kdU�"���M��6E:�ɰ��҃�s��k���PeQ\wH-{�Nv������+e �Z�ߕ����"���SfT[v�r�,_�I�޸�[L��_Xyz'�O��n}kgy��ɔ�r���.�]`0�*�f�xwV]uT1�t�"�pY0e�/ar�)��<����%�fy����[�s~��́e�D�q�fV@מּ/��&�'ېQ����i�\�	i/��x2.��O� 0���M.M̜�Y�̤]��G?9�B�ĭ)L��2~e�?�ƐA����ϸ̽{[�䶚(�RQƸ��^��^���&�@~�|"�>(Շ�tU��q��TIIK�uuu1
�ݚ?��Nn 9I�w��=��T�e��P�&ΆD��Y�j۾C�����M����GdN�d��<�I����~�!;�N)z��ͩ�8� |)�$;;� !��9_l?��F���2@��IĿ�W��*��-����2�pq3�7oor��Ͽ�w�b���	<�|Й��k+yo4~l�D N�+�����'s�������d��fy��72O(8z;�Y�e�c�S9jO�>~k-!�>x=�(��#��N}ROu����0�-��M�>�u<-R��`zn
�ɕ���"���ID(�0����v��伏���*r閦~�-���?ͭ�����ɺ�>��Kĸ�o@7�� �glC��u=	���/�����~�ڏeX�<ed�Ǟ�lwt��������g(��C)G�����ȦO���WφR����t�'�{��i�I1r���"�拽�5%F���?;�Z�[�;v?]�,�Ƶ
M2���擷{ڪJ���ɦ�GOKN�ev2��V[�,θ��[��`��%�,s��$�����m��e��KDX��9o��2[��
t��<�$cZ�j�#�����/���,�l���Z��4�(�
R(�/]V	8E`�dr�����:�N��Ν;����6e�'+����2,��ֹᎄ���F��E�\��{*�Pkfeî�'�ҍhc�Ё�K|������ʁ�ݫ��>)\�m����ӭ����rcj��N���/��9�98te�$z�j#r[.$W�X���O�&w�Z�A������Z՟�OѢ9	�ɑHEIۿ��"%,'�"˥��+�P����9�t����#|�w�JÉ��H���1˪bbbgn��.�SAŃ��\*ծr�,�I;�
���	4!s3)Ճ��������:B5!?4�Ɛ����e�z(���y)��k�ܸ�"��ar|w.����%�z_���j�#��pY���i�QC.,�;����{�&�k>�[⃈��
�e@ݫ�����Ζ͎Mb�2��e�����W+����~��z�m���/���5��1����_�s����㏚rw$��/�d ږN~z࢚�G�NOO;��Q&�����4��/g�����)�eC(Vg�PH���I�ӖN��,RI����ݎ�j��
b���/G�}+�[[۫���I*\�bb9EE���˹�*�x��� 5��>� ��*A��l�4dt����]��+rrrrdl�ΰ�2ݘΰN,a���̙b���ĹsS�r��~���G�鮩�`N |q	����]:'8\Fhu����/al؜�a-܌�� hשD<���X-�����GU����TRp�W��zL�������
�H�M��s⬣++�����Phih(UX����`��+/\.���Oϒ�?��`nE����k�ΜZ[[��W�mͼЧR�8R3�
�;�	��:k�E��6ԟT��@:�����	�[q?�����ev47W��ϑ nZ�0�1z!�at@>2��]��Ԍ���e���~�8��U�W5z.3�%/�&�F�/a5��FKڇ���e��}����ݕ�a��\�O�WF] �ڋ�l����D�M��6���"��~��V�v`�V*ɶ�@��?�P��V���\2�زL�nq7噣���~�� ֭�tnn�*g|MkT�J���+�Z�����q]�.kzvvv_��=���̡R��͞�"x����l`p��ቪ��5%̍��U����������5��g{7����4�8���E�_->tm"H��>WW���ˍ�Cw�GpE]���w��P�r�Ɵ��	V�F�y[m'����󎄽�G�SbYx!	�OB/�c�.�i�V���7����(�$������I5�� ��w�v��𳳫E�E�Ae�}����	x��Dt��\@���P=�A%��o����+�4�ɾp��t2G�
�I�rc?�鱨�����[���
�.���3��j�hv������/sj��������y�}��O5�9#�ݧ����>g��{��;J~�ִA~d��c%��hubw�l�(-�QXu6��=�0���R�8a.�)��Ш�>T�+����R3�;~4T�_扣�+�i�Ղ&�MI�R��E4M�E/z��͙�,xM_� �Z���B��}%O���j���Kr�sf�*)Sl1�z�JJJ2��U4$&�T[㄂F�~�� k�̛�b��ʄ��wc��No5|��i�M��2�x�'��?E�v�w��c�Hi������FC��_C��3�Ş$8�=؅N|��]P1]�n랏ۅ��)�+Q�>X�m�Ҙ�4������.sE��������>*"� ن�-SNmA���Ѐ��w��Aa<c6[�JI�?��U�DQDͯ��|��L�E{�F��#X�j����:^1L�h$�����N��\:��B�.+#�L~�M��쇹���G��B��!��[U#�Ug#@,��'������.J���k��F�Ƭ���ޣ[_ދ����PV�`��.�Hry�z =��+�ah��V(����4o2WWWqɻ|��:FnR�Kz��*2Y��V9�?k A#%��4_=49�0	�S� +����똮�7�퓃A;����C�I��ٯ]����m�6�2%�P�s\�#��S;Ԅ��o:݅ŧ�_k��:4%j�Tv�+9���7�^p[7R��m����{�d���%�ݓ��"��D�f���#OR�233#�@�)�x���ĺ����4�RϏ�����קꅭUR�h����E��]���)�����L��̛�o��x`��0��e���7}�[��� �C�lY�M)�����)�ؗ���Y����K���/�P��K������mԌah����S�^-(��1s�5��ԕS����]J$.N�uH~�n���T�z&�7L�^���2�Xݫe��kj�th�.ǡ�W�8ߛ�pqb���qÀP�m5:Ԏ׸P��F&�ի���`�o@������Tx�F���O���Q2����o�N衙�q�L)�����c淾o����E1
������!}���X{��m��� �K4����:��5e#��Å�.�V�0 �j�7�HƬL�K'�V�;�]*��#���m-Zaڒ�Zpu��CsQ] ��օ�cr���[m�s�u��A����56�u�<�!��cB���VO�u ��'жx�u["�Y6�o�L�o@�ͺﲒǸ^���D�ؙ�π�ey�[�!��*�;�8�W�l�}l}@a�����I&���O9.�Ҋ�:����O�"ꇻخ;�+rN����tF�׫M��Y�g��\�Oijy�q�G����`�5/����!�C�S'S!�3,��B������L��(-���w96��mP���m�-/��@��zy������<F{�0�!'�H�x鍥����5���w[�	�S-Az��6PJ�"Mqlt��&48�ܐ���F����L1�����6ވjK~o�hz�hXk�7���n�	�C1O@5�iH�fJW���;�~�Ϻ�W�Q�4��h�eKݡG��T��4i�B6�Ȩ� ���W�E��O���_�p�VUR���g(+nU�()^����ǩ=O���HJk�7<�2�7���/��@zր�2T��l���������*��4���lҨr�6M3ԛ���[x���ݣmw1#�5��;}�_�}���.��#��	�� ���:gCS���+�M���fd�<�U����9w�ˑ\W�;Ьjw�vX*��%��;��A�^�d��]�N��j�w؋��>�:?�~q�3�J@�g��bs��m�𶠲�|[>��gK�^tOtz=��nC�o��F��n�;����͂�

��6���ʧ6��3~Oo/tL��¿��?�}��ѳ{y'�#s����s��I���__�����mǧd��N�JN@�����kt�>�&QY�	�J���q83�Q��8$��l���q�,3-kp+n0Ű2��$�T��w6ss�/e`����"(�rL�ޞ��>��O��-%33x�'����u�'�ޯ�pmgq�cr�]�h!��I�w%��0�K�x��hp|Y�Q��b�VZ�~9�l�'H��,���+Ezvu���A@bs�LX6Xb��8��o����\�'�A�m�����9y�خ��o;��r�Nz�{w/�o��r���_�/�@
osn���o	l��m{��������.;�"c�: Q:;m���c^8�9EE}�ʪ;�{�Z����q-���ۭW/�=�|�s@b��N/�bo� ��_�\c@ �1~j�8�UG{�+�W�B���q/�2q�&!ッ�4�W�n��4)_�b[}K���
�!�|�qب]携�����I��dlkk+
���:� <������@��G�b�%��V�c9ʴ��Ou�C�=^�>�q�2-��!?@slq�^��0jay�]�M(B�&֪"$*t`�&�Ʀ���i»K(B�� ���R�́'�����=󯃯,�&��	��Y��X�=�������F?�u&�ʝ:]��Q�m�D
�����dee�V�) �W�6��\h��'׆*Φ�����=dw�s�knd��F[?���M����>>E��h	1����j��^ڈ�C.�.��ߡmo\������j�0�?�!�x�reV�`���Ͻ\Z�Iܵ�������W/��j�Ƞ&c�ߡċB&����@�4559qI�6��Y�#|(���C�Ҵ���H���I���jwCooo���M�w��S'#�?n=�LNN�u��\�E������sՈ��OLw��if�1I^�@i�L7�� ��^.g�ĩ,l~\���F���b��#��z%��,4s�b�8�Ք�(�c��ݬ�Z� ���C8�ם�1ʜ�\�CL�����4�7_�\&��LN�,GG'��A���m�J�\ �ـ����w�y��	�9u����?{:cVN:vqs;�R��^�l0��	�|!|������6k�}��b��\�yY[[�TZu��Zɩ4���骹a�ϭz�= ��vwNa�
,z�g�_`f����.�]��GB >]������I���ψy��Sa�i�Y��%����f��X˭��
ms�����Q`�� �Da�@/| ����Um��������c/�����ǯA "�7~9��m��$]<I�D?h�U <X�>)��>���Z�.z/sssR�J-NǛ��TX�u7�r9%g�H��^i����������Ҭ�)Ȭ4��c��(FY�r3Ӥ7�b��ڄ��^�3�`;�u����[Ho���(����ف�q��,+�aɨK�u�koW�F=��ӏ�������~�_����L=�˃���#".�O ������%j�s��ϩ�6,���xE��6u�U�@�ǧk�����L�O�S�EY��$,�I����8��S6���"���w.������'My�&��}���쭸�o^�!!%&��5���t�rf�7Zi?��~�̩e7\�4X��S�c�.��뵐I�{�L���@�u Q��`�O�r�VۂEM�����y%ۮXp�;#��	g��&��/Wy޴%��ɻ�,A�1RB����������<��X��R�?���/7�
@�/������s���ڠ=�7HHHH�����T8[�N�0�P�bqN7�(�MsmT�<������E�74�a�'+/_f/����,_!�,dDP'�L �\v3���݋�{��ak�_��]�KkRث��ɂ�u��I!�_�.�fی,�%n�W��f�t�������(}�Bi��^�
��z�ʕ���t	X���?(�L8t촆sx�6�[���p���gQ�������"�>>>��ɐW�����
$�������h[ڡ�0dDJf��<wf��+6��#o�������ʍw����ƨ��۸c!¥җ`t��9o���4eL�Zm�dQ
͐r�չ�/�?agg�(d|�1U�[i��8��0���VW�]k�HL�/X�<�031��O�"�4���Z�#LF�c-��Ɍ�g1A��p:W��E����}���
�k����Tq��<-_i26��&�%�?�:�U��#QL���7>p,C�֤Bv�=��!^�����H����#b�r�I �'��E��ښ�?��M�I�v�ڿM�@�N�)�����[�DB��YT��mLY�X}�R�zg����� xpp����wfo�=�K��ȫ��M�".��#`�^?��t�=��>7[���d>�Z�/����\�F��k��%�I�̜��T�����l�V�����CG�� �Z�-�V�����Vw�h-�z�BX��{�TG[[�A�=�WX���O���d$�����"3`�a��Tw�jx2D����A�er;1�B�W������j�j�����4i���h�H�`���ٔ�WG�-��~�e�)`���i������������6Ѝ��1;�CC��PK�p���稝~Y����H" }�A:;D�E���8Ĕ�`�n�we�r��*u[W%�e���6��χ�ɢ%��u���t15��Qfԭ10�k��c�򻩞��} �+� ɪ|�A�q�5A#�V��I�M�U,4 �hg�"�ѭ��{Y1���F`y��:&k.��so�N�&᳡g�����6K:`o}y] S�dJܶ-�)p{K�c������"����-c�@:��4�ukٷ�]_�3ݫ��� rr��B䡂W/P���1��7�fa����:��{��f����z OM�ю���Ke��O:��}�DY9X�#�8��5z�b�׹���F�@zlp-A�0�!�os��6��]�iFF���j���P	��ϵHڝ�w_�6��ƹ�A�%B@eZxznsr�����P�|�-��D��d���ә��)��p�����e��N�{�UL� =j�H�� ����I��Ƽ�����;�Y� WdSǞhR�J��ߕ����ЋC�� ������Z�:�5c>� �OUb7�6[XG�(6������n���$��6�����Q��9_�\�}ӯ��K��F�~O���l�[B�J�\VШF�Mʕ�:?�=�_<1�@��"g�rR!w�X�&A���!;��er���L��]}�'"-"��<,� ����S�h>,�R�TnBe�l�G���TCH�U\�O�!�m���ɔb34:�J4��zi�@:X�PgJ{_�f��Z��聼�d�7�Wm��.4���P}��u$mL/��� AP���g��,���)�A'{\���x�i\A�~����aVi�x�>���W��r����	��kȿ0��Ł�C���35��7��9���=
"�~M����[���b�O�qC�c Ĥɷ��џt.&#���=���[�!����!��6뉑?�w��:�b�4[�.G:'����OCo�*~{Ѳr�������&�q��e^���l���/�^��f��
.�{j�j�]���ͬ�s�w���7��sl��Lȅ-90�+�� :�ݳH,9�̠����̰Ok��J�g��-�	�ջ�Uj'��>�dCw��u�9���.��Ѿ�؍-f5\l-Lybf�HȐ����q-�N#ܙ'4�eת��=��Q���<����ʌ�%���3�&�p]�ר�t/��D`4 �EQl�:�+ah��T0,6�L�úuq���b
�7^�aֶM߻9k=:�G ��
����4�_�pqvg��Dn���n��� V�����w��zL. #q��n_�޴q�mQ������ n���_�&/��
�;�ZA�'���@�u�{�;1�~�փ��ա��͡<�c�l�S�M�����������D����l(�s����|���=u�~	�dh`�X�q`�}��r�������Oޙ ��jo�B�VỎ�&�/?��~�_��+�+��T8Z�4X?�*��oO��\�W�ڄb�yO�pɧ,˅0ˬé��rVєh�dI g1Q����E���Nw�ɴ��q�!�b���1�o({;=]�i�p/��@�����}5��K���)t�H�M���X�q�a=�W�k��*��R�c��&3�cRB�|���vz����� =�ȿù��(����'�I�sʅFp�J�"��;���n�?�Y&�2�4
F�:��@l;4��g����2����c1�������N�	:���~£�{��R~���"_ܸ$<�!���k*i#ccl̖�rQ�+R�<5?�j��S�J��Ɂ��nmlll���8W����b�3��̈�� ��$�����6���E׊�]�n�(��Z����*�u�VVV��9�<-�Xc�Q���hJ�^�9��P�MMuu��7��t,aã����zS�5\�S���
OI�`EiT�����8��n=����v˭��2-D�ȧ�-�lSm���;��Ƣ[�T�A���ձ��B)��K{��X���ho�x�U	�����1��T��L�"0�Ƥ���1�c��5���4�\����`YR��ꫲ�`�T���Lg��u{�ܾ}�Igg�|_|n�'���Mپjmwu�Xoh�I6x�+��l�q���'����~&�<���x������e�aU�Xଢ]�;)����t����={���°���[�T���*2���6��z�ӓ��Z�5���0��;�|�_��������ÃA~���F��)vs���P��û��E��@�s��Ff .�Yϥ�y�
|~�(ܰ�D␡r4���	'�+s��Z!!!�T�����Y�i&UV!�~/+w ���~M��X�?�VY�Ū���> p7Ӻ��g�h���^�*c�&�8�^�#�<�@(}���<�:8��qw���{����;����c���5Uk�zؕ�GK��h��q*�JJJ��b���Y�n�3��E���z��q>'���w/�8o�%�I��֔���c��؞������u���l�Ԗ�gq�"llY�L	�����8��ͤѻ[㯣����PE���,u�1�����
;�qײ��y�����k����k��Սmƛ�h�Y�V*ܭv���i�]�sق9�t�j�Տ�Ed=����ק����5kRL+(��c��#gf��`0\iG���̹)��}w''��Ѐ�;w��@��i�2�9k���� q�i�U�R���i��M�����z@��mw5`?wƹ���N�g�m1m9Ʃ�����#��=�L��3B�@ Z:����㯂ӓ,��I���ϝ��/Q3Q�P}�E�������3F4�)WR���)�b�T?h]�}'��,μ�|!�,��s�OZ0vr2*3$0pjoP����k���(�th�#�x��M]O�a���	Ĉv��@��U�E"�5�	�;�\��{��ϫ����*]�SX�� b	�7L]�}��|�옶6��ߊ��G&�nS��bBE۾��4�b`2��O�{�g�xRF��s��>d��/=\��Bt���������Kuyy�~�M#]���m�ֽ^��<�e�Z��G�k!z����X]�x����k�Z=���/o]:��;�����2�&,l�?���vX�[���$n����k ũ�ȣ�)�Ȯ�o���ozۍ?k���Mb+�z���~�ӧe7�ڠ�-����C��3�Anj����d�\�oۜ��������ex�J%�J��1Š�>-/b���P�BfWa�����k,��I_6�H�dm~���3��h:ؑ1����������]�o�l��Z���vL�ɌH�q���RI���jvt�Gb�UQ
:���r��j����@`��w����x������=�2������w0��ak�䯼H?��g:��1�.�ߏ ��H
��w��ι���q�Ʃ|�c��U_*���K��[�4&;q�q�Ht���8�E��e�~u�bޚR�tQ���,,!���(�T�����J��);��1uy��R�xw�tM���v��\.�	�۬1�2j1�9�!��uى��@�4
��|̴��c���m���"Ը.�ʺT4������5_׿N�=r* >�N�.Uo"�s���p�'�}Y$i�� �-P�z�Q�ɘw?��$��*p�:�=�V�X��˕�/�䂒v-���rF���E}�f��e=�.��2٬�5�۾�=i.�^����;�Y��*�ܝ�)�z+��N6�d*><���2/=��E��3��r��K�=���@C��sKEn�w<�@���|xv��B_wz�Аs)����~d+E��\c�NC$��Q�Ob9Fgg��}�5@���LQ.z-���=F���%�6@��.������' ���ħ���yղ림�]~TF|�uG��h�_���
�8fn�҈����<kϧI@�}���P��y]��G�<�Z7uo�U���ʩ5Q!��pj�s���;�]��]]���N�|nS�ͭ<P^Y��*0ЄG3sd�`|۱@:�<_��X,=ϑ�{Ӓڪj�|�z�����Qf�ｽ��.�/B�$!�໅������Ik#�Ad<LSA�o#]�`0ֶo�:�,P��7�'Tv)Q��9�x����^Ӳ�����,Pv�*Uݐ�LM�m=4v�6�_���z��Z��SV�N���K3��B �dB��zF.Μ!�rĦ�{�⟫܊c���m�(l��ˬ�R��y��_�U������1^x�`�3#ߞ
��K�Y��pg?�	��}��~�Q�1�8#BKyl�n�s�6�HͲ�̓�A���j�>Vb�����_�����mxD�p�ȿ�Lu�m�������Ͱ���e��}���a%]�Y����Y��ѧ����9��ˑO�vs�=Z7�btv÷c~˚�U����m�J'���=����?� �W�e�p����b�8s*t!Fj�G�G��&=b�&�S8z��t�Z\��@�ulku�N���^�K����:dܻ�;O�U�h��l��Vʀ��8�v��w��	��+.7�CCD��|yDj?�;��A�[�rx�<���	:�M�I�{��&����55_��$�,l{{���9D����a	cv�;)Qc���>��`���̳f���c�m�!}Z���r�����g���z^�tci�6m,��w�!��/|{�(��e��r`+ʴ.}��s[y#��|���\&=��{���a�1�j{���_h�74�^����mr�Kni�+h���J�X��'����>�ޥ0ĭy+�r=�4�i�{����E����T���?�6�'�3I�����.������=�Z���+����NE�s�Tt����Ѷ�W�k���#��t@�/K楣�TA��\�5�]��5'�T	_p�0������E��O_�-�2�{�O���xW������	�=r�Q��^�&��N��P�٨��`=�`����S
MGoձ�%�n1n�X�12��N_Ɏ�<�
r%My�~����r<�1M�X�Ǘ"�8p��1�__�ђ�����}vo ��^�q�LT����g��Mj�o��	��Hx|�/r���1�������Ze�:$RC�����`�|х�vnL�q&�I�\�w��,��=��~u]2����P��M��"�XV���@4)E#��uz�:v�
h�#�-����&�(�a��(i�1�3�t�hq��@YYbRy 7���np���1]�؇ǋ��|\]u �����	�,8Yi1��/���7����z"�Pc��j��X��.�~�8�!p���Mll�]���t)C�7����X��#���Zb�I�'kѢ�=�R3�Q�/���.]�����u�Gйq��bj@�c����o�xe�s��2D�Hӫ�P�f�%�d�����?���*K�����������yE���xdk��ƐC��(A�>�o!�(O3��"�X����s�ǌ��Q��X��ZF��9)靬u�����vk�ϟ	�Q����z���[�����,08Vj\:�k&?�r���a�Fò��o����y�i�k���h#��	~�222U�l�u��ճ�!��Kinw	8�8k�C�������~K���*�U��c�c�w��g�2��񭏟l�	rϟ
5���~beg{:�Q�V������aT(��t�^�[���	~� ���S~���]�9� �q�_@] �%i�*�O��]29-_��t�ׇ��]��x&�%Û>׆��dvY_�	�����Tt��+�U���v�e�]������&fR�Q������|q�iӶtt�>�C�Q��fi����!�����������:s|DrZ��0�YB�8a�$	u)��ֺ�����Z�X�3ۤ{ ��N�|�,iK�C�]��6�T���5�����D	��ѭ8ol������:~'�)����<ޔ�V���L~�]d�=�����X��	T���ݨ���v��a�'/��w79�m_K����17ooݜ�8��!nņ�9�铎�0ԅu�_״�*�N{�O+v`��@}�2�u�~�Lȿ��A��ԣrf:q�w[g ��̱i)�!A�
3[�O����w/fgy �BU�J��a�ࠟ4l�`j:$}���������G��ܧ��0m�������R��a�u�f .��n���mx>V�L3hM4��\F[�ӧO�6x-ۖڹ���=6�R�*�j�66����Ω�φ���jAS~?���Q.��Ւ��=������_�
�kE#X�l1�������T[�����ha��U!��;p�v+c3�N�e�N����}sl2h���g�����wz}��#'�Vt߭�=��.�̓X螁a�W��{��c�������=��d�tx6��� ��8TN�o4L-,�ZT�6-{�u.����u�ӱE	�.�H�����]/���<�x��͋�Jv�R�]�6���^O9�#�[���*��9Ga���ᕆ�{1�r��2��T5���B�^�������L���Ү9��vt쀻��`�CvK����#�:?\�?���x�N��{@��`�y@��f<�wTҝį�����w�Y.S�t��\�n�]�*I�!�!EDx�$��1�>�,fן{��`bT똔[�5�;"��،� t��.���HqyKj�L� �w���1X�:O��ƍ:����vY[?�!j�8��	/
�Z�wQ���h�߲����g�q����D��jLfg�_n��0[KO��-�82<�X�%V����8Tn��@Ny�5F�����O����|���x��"�0dmn�x�ʕ����"��p�A�Q����X>�#o}��
�k�hh7������75K�oP�X\�<K�拦ځw��f�����6
�'?Vm5X�,�g|��Ɔ06��.n*���Zf6��U)8�5F��E�,�9��l�EY��Pk�J\X m��������#�rӐ�x��z���'u�2���� �� �� �U����N���!��H^14S��:��3�}��'d2y�Z5�L�6����� ΃�����B�CP����c��𔑃��޶�; 3�Uҷw���k�C���rr&��W�
�r���d]Ȃ��vk��-�
6*oގ�🥚���ؠ��4555>�D��5��b�����!Y&`��a�{������ŷ ����B�ϲL͗t�I�(y�Mܱ�Y�{��﹠26O��5���Ay�!PN��Kxvlȟ�UaO��l��y��m;����M���e�װI��8���_p���5���?�TH���qCFk�"�ֵo4�b�H�j�����mo7Wn��z���2�}�}�F��:���r��c4k�*���h�����lׯ�d�f-����Nd8��%�A����Xu4����VUՏ���������r4`���M��1^0X�J����UaD�c��Ն]ݽs��]�f@��z���C�@e�zQo�p!�����
�y=���^���4��.���Ӝ*��t󎱻�# �:�2�Zw�H 3뀗���ZO���D������.�Υo2����^�yc��_Iy'S��{��j�9w���@)+j��D��M�Q�Ϲ���J#�S�^^�Ą�C�u(�]\��*��} ��pJ��������0��ժw�3��I+��ǳ��ë�6�/���bk2��(�w�Z�K�6�hjj;�y�.�}nʣw C� �Fk�~ʳ3���28@" ����2Y����Y��QyRڙ))�?���͠�;�� ޓo�ws8�>��˛?���-��Tm=;�����g�V�N� ��o��BT���UK�?P�v�0.	�z����7鉹��j�����P�J�=�=yC7˯��+���^ͷ�6�_R�����q�D�Ծ��JJCf�򏚿֦���]�8���u�GP�X0��+1������c�p��FF�ㅅ���$�7]� �6�r�c牧/2���Z��P��t?\6�띳�����ÿ)))M�8��~vEC�P�/���;�f�P������]�/;)N�W�E�Z�: ���oǮ�����y��:U�(�{�G#7�g9�w�o�)�v�m���c5}����b2ߜ8��{|��p�\����r����D��G���֯Ʃ|ۃ�|6\��a��UT��*\����_�m��i�R�^�M)Y�E�m?�r�h�}�=�@2�j~����Cݏ��KF�,x��"�0�jv�n��:�8vr�{�&�a�!�Q���筭�x��	P�qq������)q�~0$X�Т�����)�m���u��5.��O��zV�ֆ@��._ה�z����ӂ�1���ʇKGKˇbbb^-f����@[�m;��}y�r���5A�z�ŋt���%i7������!�RN�w(���悖 &�m�1��fì�HeZQ9^�i�zT�DN�J�:�gü �:�lȯ_6#���"r����������y�2��#�tNsu5�@@y6MGu�7z��3:����WR���>ܻ�Rg@��S�n����"�=�Ψ�6frrr���͚N��sc�4�'O(�G����ثb΀�°L��m�U��{�L���0�Jj^��6J9�}��Poz0.}���yP�צY�,�A{H%�\16���;��=�����t�X�L�u�BNmeO{��~�V�	z��}'���Ҳ��I*\ޫCy�w�M��.l�� ����>Ce暠���?�a-&��N��m�w� +�����8=,��t9�oЊ����<��b����[ILT��>T��-5��=�Zލyb�C��Yj��*g�9�w�����>�#/�L�ۣn�}�ǵ�鯿|�<��	:ժ�����N�a�����h렙\8!-���������޴L=�?��k{��՘`����*�\8E]��N�M��hI�I\Yp��S�U�7�1ŀ�^��z6<��
0���lL���09�\�`h?����ivy�t4�#��-}=��]����tF�dx��]d�`��S%�aJAF��~�o�+�S,���"�2��Z�/#.��i�b@a<>�n�*�pz � �*6YVF��2>|N�EE�������;h?�O5ܕD"ّ�22|��CҮ��NHH�Yqtw>�G�q �ذ�ϣ[�I���o�^�V+����ޛ��������υ��4@k�XZ�H�dF9�G_��L��fsk�M�x���Vͱ��AW�(K]>�m�<���u9JPP��A�E�S�MbD���L�|��͊uM�;�IG	����Q9��Ie��+�Ism��wWp�}%�2�x��7���A�ǀ��<Vq���;�6R���M�x�+W��W��X�n�7n��<�Z�_�`�� 	-�隨����/�&���V�?!<�{{k�Ʈ����$8,�3����[�З��U�R���M����A��9�<]��b�>3wy��|�G,x�UQ��Ҋ`2<C��ts�=�g�O��+&�k����My�t�ZS�c�Ԙ���H�,�֍��wu}\��
�<�9�c?8��x�N��Ud�W���^<����r�7�����XÀ�'�0�ص�0jW�y��9>���p(�d��>!������*���9 �����޶��L�-�����QH�����`�����>Xe����
�����	Q�RDI�P�%DZ��A�C�����n���!D�!%��;��}�7k�r-����}�~������n�ngf�SRRZ�avT�MG7�"�?�_���J!F�����~׫Q��֧³��e�Q&'���N!嚞N.d�l�m�Cy�[(���h��ִ�S����/�`
>tG�����S0'���v����;@kg���¡�W��%~9у������j����tu�菇Bӓᵒ���#+<�����g	ZVM�]�JDDD�� 7��^����<����+N���l����e���{��1]�#q�!�����g�"��6rBw�$ U��I���w~u����i���~����b�pgqͺ���9�BO�ָޘ
jS��Poџ�2�n3�ZE���Ɔ>�����g�}5*�2���]L\f�������#ex25^޹>H��C�>Qv��1#=]�t�<�~�5'��h~� �o��d�q��n�w:[�yoK�d�8+�9����e���a�;�۰����T��[Cf��/6��&�L9I��Ϣ����)�{�((A��B}q&���H>X�7�����nf}PO��W��m����^0,-ѯ`��X���ͧ�#��;�������󬓏���i��H�LήV46�>�t}�<�mk�ph[��[�Pi�{v�:�hk�v�h��D�G�g?G��;���s�riy�ՠ�ƽǻ4�o:��8��$�����wG�����d�h�+ZS����	fk��Wے�Z��&2�}� <<|o[���'nQT��ϳV��Px��r-2h�:�E�\�X��i/��ܗ�7�*��P�q�/,NKK+�9�3�n��O�q��2ŊD����gc�%6P���UWS�}_� �,�����6��g��`Jk��K��Ӏ���Y����:�3��<P�\Ec_Lk0^���֍�J'*)sU��+��uu�w%�VY�&(���Q�,�H�������FNx~����������G�Ĩj4KH���H𣐣���4���3��ZR��R�`��o��Gz�/gr�?w���(�}p��3N����V|�
dyHG\��S?	 bC�RKlA$����B���By
�읜�dV�[�7x�Z�'�ZSݾ���;n�	����rJ���l�܇\��ٖ�9��t��~��*�Ç��y�j�8�Y�L[(��Im�6tX����$a��ڒ'
�W�d����LM�׸�ţ����ty�.SS
�yS��)cri�=}����`�b�Qe�ܜ�NN7v<~�%f9�����RSS������.�i_M:"\�c�ż$��N�SE=yЯ�,hY_�����ayy�(z��d�.�YI�ޘKTW�`�R�5��Ċ�����Ф������ +kk��m��'w�
��?�?Ff�����dGs��p/;��f4��5T��-���g�/���dб�;j��̴K<�Χ��<�2�ž�:�Ӕ�!�U��!V$�tr7T7jPj������N�v�z5_m�{�ߝ���a0��~�g�fo����vT=�3}����p�Ս�G�gN����������S��&�����Ʊ���Rs����*�e��U�N���?�H���y���ǼӴ�"Q��<�y��@J�� ���kŪ��ď��+ͨ�ǉZZ��'wp�������K�W�-�,����&����Z_= ��=+��N�(�g�W�r��� S�]t�DHWh��p0�/�àq烙��<r��L�`.S��l�e�������~��X������+]���@J�S%�n��9��^���Te�d�Xuߧ%��<9D-C7�2V�|�R�	�7Չ����ƺ0��2qBm�K!ɚ���MƵt��T+�9X$�Z{.�2U9���b��6a�����w�:M{��g5q�h��Ɉ�kI?�ᐭ���J��y� ����xKK��6c��|v� �j�t�L��Ht�;V�}��=ٰ̼;`
�g����3��(bRRk�C]�l$�@�}��e�����5��߾ٜt����,'��89��K&��NFF6ʙ�m~EP�-�nR�Pcj]�����c���s��햖��G�^�����V��/Λ?I��Mbyo.��`ن&h�4ӝ̬oP����>�.��J_b���)��'���q����F�^+!q~�xD@�'}�N�{��q��q���Z �Ǵ�L�x��<���37�}���1�ʨ���R��Cx�� ���b�G�a��#ūR����127u��`y//Z�E@�������D=��R��dp����8��Y���bɵk�9�+>�t��B܀����]���=Ewxyߵ��$��~;�� �/�հ��k>�5<����=c[`����h�iB r��刣(M���l������4�u��[4c�\�����Sh�9�8��;cWg�r>�X@'!8/���z���08A>�}�'�Hqҁd���ۄݹ	��H�m^�����npn��G�����ߨk���ܼ�.�[��^�@T7�S�T�o�57/��9�h^�!�OtY��7��fη83]�R��YW�t���g��,;џ7�i�*'{3k�?�,��O�]��7vqF�C��K�k^�/�֪BA""~)A��hp�QH�3�!s�Ϲ�aU)α�W�ZZ�
I/{����ÒC������cz	����+.����?�'�ur���5��� ��*++)�0�ͱ�ٛ�:R�����(��_O3=ٟX�����
�PE��JA/u������Nm���{F�ӱNd�fzd��`������(|���`F�\ܗ�@o`A��"�Wc�����'0ҁ�d��bP�Y�d��&O�F.�t~(O�p^�IiJ��>�ce��RZKK�H���������ҁ�s|�]�Դz�����K�_�p��d����v���y4wZ4弛�a����u��H��DﴇE������B0���J-��i�Sm|E��E��EC�td�������.o�P��[����|�NBd	<>��Ť��_�����w�;(j�P��b�T���'�����K��r/�ή��Ti��`.G@��K�Pm4�7�����Yy��r��͎���-�; ��C�М���oHEOan�wt�]�n�������ޞ�(�T�+����j���j%(U�N�t�����|zEO�>�w�Ա*���@+N�k*Z�\�u-d}�M�O��Iȵ���cDk\�c�!!!�$-�QM���ͺ�fݲ@4|�VXh;vV���:�����h�r�A�_��>�c�/S������E<�����W*H$���ՕR��q�i�1��^�����>wq����2�6��Hi��� sA�-��o�i�|����x���X�ڵ��dWU�z�0���ӧ{�]~���� ��}HWe�-`�r�"h�I�m��E���@j��Lt��*���hC��3:B�gn�J���࿰���� as�qy��2���Ʀ�+K�$ڶ��y\�vk�h��LYx�?����L���e��VNlI*ϻT.�k�չ�X�~��)�~"��Q���!�����?t=��X�-�pV���U�2 ����tX�*��2��<�ֶlx���[q� �M{���{����	��٣?�����`5y�r�������;�j?��<�(,럙��>�k���������g+�F�@�s���@����i�5b/�Ve1WxTace�^���=��C�3mCS܏�$��hי-�D��;�vff���_9�9�I���LC�	Iע�N�2�!��S'����.��D�)E�pƹ�M�P	]0�?�TV4�i���Ⱦw�Eє?
��W���ev���L�);z�a������T��=�^���rmP��/b�d���X\UJ���Q��MP�^K�B���/�%���XMkU|�n9{!������)�W܃v$Y�~1��=C�8����]�o�����!���֔Nđx͡z�n|s��@e�����*��>Ӎ�o%3�N>�E���8J
k5�^��Xu���"m7F�ihp���;�V4����`��mv*o�����ʋ�4-�^��!P�C��=Y[���������g�}"D�Q7���9'�\Ӿϥabv����I킧_4Y�a�&�w��3�G�� v3�
��i]�/���O:yb�`�l߲�}�+N���TWW�PBI���<0��y|3;��B�V��9��[�1���t�_���RN	NO��<�2��1(u�l���܏��\Y��n�fƣ3�elb�H��>Hñ�Ib	�v�t�Gg~��$�Q��cccq�o%�)��$��%�]��Dc4�O]#xp%��7�fg�uj3��z����՘���-��	���d��ɚ�
E V@d����O�ӛ�6*2�Yn�)��ܿQn�Ay�0&Ӻ���x'�i�]q�w�(Xұ�(���$3��ޭ�ԁԺw�C�������F��QK�_��'�x���+]]2"�`�:e��g�ISVpx���G��t9ơ�I0��ǖ-̠�GJ(V��Y{��	�D�ǨJ�{���x̃7�Ē��{y�|D�x	�Xc�I(�`���Zce�ȵ� �/�NӅ4�+����Uȹ~w0
�3�tF|���s��~��������l֕X6�z������RG��JY�����O����������>~-7/oxv�c$Ϧ��9X��g��Rd�R�־�wV�YLz�-��ڈu��]�P��_��2M�{������l�5�M�c�Y�7��!@3OO��^Rj4�`O�1��v,X���������d�$���?nU�t�spX��a>�C�Wߢl���O��?�β��A�gw~��d�� ��9����uT��٨�2�ǩ��nX��F�*c��N���[�jg��_ڿ�;� ]6�?Hf�'ѣ�S�8-3�!t����j�ޮc����mL0db����iؒ?�tr��V{V&���-�9U��8�N�
�I�i�ɓv�k?ϴ� ��B�]�X�ۆEB���!��4��������W ��<өlsvB����x��'���I�՜�����cDC|�`���{��߂�Ju6�c徴/�^}2��յxѵ��otV�sh�TBz7},���i�%$�;����Kh��2�b�<���D�WUV�Y֢m�2`��gf<,?i�;4���E3 �֣�C4d��c�����"k)�=)�L���eR*F7ظT���p�Q��<�|��l�i� �?^��
.�κ��m��~f�w����c�":���E���{s�l9.]�;W��5'R��bv��{�CҨL%����2?��A�@�j@uۮ9��2�������h��57K<b`b9�Z}Uf�!D���KTzz�{���U��p��|�
�O j�>��`��`����f����-W�E�zq�S)�J�.�˩�ƶЏF�#�����or� R�c�]�)�t�\
�^��ǃ���O����~�-7����'wl
�p������v%�{Ic�W�	6+�z�%���,����˰ڵ�6V�?z��)Ò��M�m�7P2	�+����]JRR#FR��)�$7^��g�K'E�
��������#L��+�<>"��s������f\7�Z XB�p\��+��u�ӖC�}��qRL}�����*�y��aV�<��|cTc_1��3����1ȥ�OB~\����cU�ez���R1���Z͌�=�g:�^��=���F4I-+퐜��P�`|���M����T���k/�Gx����}X��0�͈�����6�|��Jo��U�y� >f�,�1cW�ݎ���j��E@��u{)���䢠{n�	:���۳5oqܕ����3:�F�w�8�S,ε�M�٪9�dr���
�|2ӹE�����/ȥ���`�������I�Kr�o�BYB�X�[��N�MnT1)5���^ �w6v��ˋ���	)AK�7�{���v�븧�k��'雺�hJ�d�d ����?�p0�;�-����8��[G�;�U�L�q�#�l|]f:!���͆����d3�{���*��E9$��{ׂAN��	��o�{j�X�]��b&o��s�@�	�x`���j-#�k�yy{�]�u<=|��j<%����茢ޙq�w#\�sb�}���z��� �1��͎��ؾ���丫�����ٗ��.��U=�ʚ݁� U٢hm�Gd�,8~ll
A%�����6��y,��hJ+ �n3��hX�ﴤ��I�D�s����t�G53<?��h�8����S����� 	W�a��Rj��������߷�QC�0J=Vu�E����řŧC}�2A��h���rQs0e�z�<q!�)�%�.�l��k۱1>��T�ےhΜ�fzA��M��9F옮 �LE�[p>���2�5�����D��D�;<��n@x%5]RO"&&v%�0����aٝ)�ҫ��@q�J�-y���y��;�f�J�ޑs�EE��N����q}����#��W���
$���g�j����Z(�!	�^@*F�[�!�Ǵ-����F���!ٔ$4�Ͻ������}�xY{��9}�����{GP�G;
م�:����-�,8�"D�ݭ��`f�Ieddc2ܻ��π� �~���}1��f��~���I:��S�)�&��z~��urH�7�WA^�������⻷}�~������"3���'XR�)�>Q�C*�SN����ԛ�]ZZ��vP۹��9��&�6P>N�#hJ-o�x���?����d��'�PKc��VNo���C�.�8����q�o��u���|��h{Z�\#O�U�'��{�G�y�p����[y�z�z�|�hG�]R6)�4_ͺ��,�4���u-�b�B�>��x�_�q�5:6Q��E[��p).��УEN���1M@�p���Zz�ٸED"�Y�+D�Ed���z�Y��D�3���L����p���'^���N]ߚ˯��9�+�4֣�}���S[.��h����p����z�G���B��--0||��1�����瞩�c:��t@����}}�(C#�E���3<�����.��Kc��8^�	��	f�dD$�5�M<��/�� �:Y� R#
��q�r���8�y�F���.8
5�-8uDP@;��G!!��ru*����4��z���b

X�HH����տӱlu�^�7�@����?��W�+hիq�^������"N�:+��}�=.��/Sj�/�æ�ҪoZ�R�~#��P�N����$F6L�,D#I�i��sݭ~U��j�<�|?���v�*��h���)x1X���%à�+я|���N��|�ĉC n��f�?���4E�q�>�W��7�P{WN��Hh��0z�7�
�)�噏��ke+m��c�_sa��C_�[M2n�ϳ]�qV���O)E`��d�}8[�"`߶ܟ�z-'���0���X ��|�F�����a���b	��AM�T44߫��6�L�v��K���O�o�� �]����;E���(-C_�����,�Ñ<�` �����V����P]��r���}�@��mc*��(,���971���}��Q-�hښլH 7���}h�]�^���(ٵ8�v"�m�vI8؈Ђ��;&M����P}-x��%5���q�e��3��5S�n>�R�_�d`��loI��O�$�Xz�Ϭ�P腍zL�̅�=�?�#�ek�fX|t_����tY|�?���;�n�𧗣�3�/���L����a3_�L8Vj��or{�Җ�m}B5V��~���;�~�i�E��J��/0��-��Ք�y7��i�����P�K�hu��
>�N�pM�����p\�	{v�ѥ]�1b!i�݁���l���ki>�m��oz�xUp����2���5v�$��<���/�ǊuCuj�olLc��#�b��0F^^w|}}{��F�u 0�P�.�K(���P>.�L�0�QA\=�H�yz��,Ab�c��Y>+z؎J�� ��z	22nG�l�M�8�xw�E$���u�(�>�?�5E0�u��!#K��h�Zws���Z�z�MQU��<�}�"�2l���,�r��:�ik"]�{;��(C����/�V ��hUV�PZբ��h�\�g^������v��g���Z^�RoQ�.�^�����{�
�a��&��OW�$v-��z� ��!
\L'{zP��'�{�v�kP����F�_�����Ѡ� b��5�p=:�+�{)s�˂5��;��,NZfP�6C��ݱL�{��q!�m����/44�nY�F��m�����pN�gW�ݼ5����Aj�(�D�F0�Th`Z��Q��Z#�p� �:��IaN��K��g�L�$�tw�C�f�]�-��{aKx�d���]�p���b��������iR=}O������qǝʔ㓯q��>�b�?�����n����>��˧����;B��o��{��8�j�4nu��>�����po�=�pq�c�1_oX�]�G�_yN����V�:��@���k��}1(�4{�B��޲��#�,F�M�N�w��<�^Ų7A���r��ݺ�>�˓��?NӅ�uwl�:I���
l/���WmC*[;�n1,e�O����I{0}3�����;�V��j�
�<I䈋~���y/����*��@�x\��2m��\�2m�C\&4��Bi��&e�8�I���=��Լ��Tc������1�9����� m�B�r;��:�3/�T$���!6_��o@j��Agޔ;�R
rr�lǊ�%���,�mj��قww�<����q�E`��)�pۓ���E�����x}#6���Z���2�Zi�\!�z�X��ߖe��p�;x���T�)OB������:�^΄�S�0$�IW����yt9�+ ����p���Tr?�,��m:Ӱ�]�����RR�c�Zmb��;Bv](^����y���5��7�*a�A����m	��I{���C@x-�ny�n��1.�ý��g�滙2���AvB
n1���KIZ�/b��-�̿���+�3�F��gUT��8Tg�������qF"u���˕jk�d����:��C���^s���p�M��5QV|���n\�4-�5�o�EXi��f"b����)�Į5>T2"�	[�f���%ᾩ��A>sM�E�R�KCCC�� �/]�51�,�互k�p��ǻR��;w�_���ar%XRG�_�����
���;X�oZ�8�������x㯅hjE�$��B�������-|q���"�Tk\�9G-.Dr��[�6Q�ٲ1�L�O� �1?�)-m<��Ѹ��[eeNPw$gUcN�ݿ'gC�PS��?����6�$��q� R����ԅ�tq]�3Ur������z���������!V�����+7K�}3���!���B��y*dv}x.���e)����ǀ]�l~�s�M{o�k.�\�W_�^74�q�}�2�{ute7-B&[&,��P��e� PZ���ճ'Jf|n�������������~DוD~S�:Ƴa��J9k��<'��x�K�U�q����iZU�p3�w�AP�� ��V����܅���~��1��qAR�`��ں�AEFp�E{�i��(�2�V�"�
�z��΁��X0`�V%A���֧>'�s�1%������>�j��_�Op���z�/C�y���� ?t��22��lv�;1k�=���5�"؆���sE�-l/��	J���B�Mm��B=h	_��-D]� �`��=y�����(^᪒�b�ڧr�=���"C!9圗u��f��SJNO�a�W��C"�c���	��u+��Y���GL�Q�.F�&9���F�;{�T�����+T��0�p����!K���H\�6�eu��?	톥�=�I�L{=��C�]>�FP��Z�^}���k��!�&%~�Z���'"���� �,�&��	a �u�����$�^�/ ���lek���F���&��[z�;(��Q��H��CǼ�d�h%C�u�]��F+�[@��R����6�f�:4�J�ZSgO�ҋ��>�"k�ػ�k�����L������|+���I�����666�[Ck�=�<h�������H��@H���}w�2�mq���\3�n�]k��	,��:��ZtB�Lv�V�	�}�u��v<h$��c�N������6�y"pH�� �{�ȡT��]x���I3�WW������i���[�Ϸ	��AMؖgwFGG��u�-����lDh*���)�B�7Z#����a��?]�Uz�J
�J,I�:L���3���	o��ܾ�2G���>�p������/?�>n �4댭�@-O\?�+<,�L��Tʅz��q%t�v��3�ϰD�sE�p=�._'���3�Nh9P�P��e��[���<<��w���v�7$'�oD L@ ~����9���>�w�r�4���h���,cL��HY �cWXiHڷ0��tv35d7o��=y"5:A����rv� ��WHU�d�E�
F���,g疢~�g�ڃ�^�>�>C>?:)�$)�,�����U��QɅ@���@����^������s�_��gk0�i@`���{�콃���Sw��`-ت0��Ď�|\��ϟm-�!ˬ��1��%�-�s'�4�?ӑ��l���
b��:3 �_Ϡ��~SK:����}\���ۥ�m�`e��A ��.nn��jir�ۿ?� �kYs˷����Pݎ���.�	���!$R-;�1��!�l����9��g=��RI#��'�ÖA���i :/�O>R�ż���4�]#g'� �4�g������=��U����Uڠy B�&���LCVW���������n��q^ĭ>����`�x^j�xVΞ]_O�jt�Ո~tx(�66P��
������1�`H��� ����Cr��*i4��5�!��i�ḃ�e���xucc0�+�؞�(���l*Zڴ�Y���5�6�~ۂ�H43U(������ �O�ٍG�a+����:])%��=�oUU-:�����߄��eZ=���5 ڌ'\��4��F&�k6�:<��L6a' �B4$!��7�^�O�J��ᆶ{GX$��T�Q5��AMRY2��p���+�z.�5^��[��^ؿ�����o���+�_��/إi�{e]����:�?��b����F�����#�wG��VLr��6�h�8�L�a�����	�l��� IuƟ_޴���ߍ��KE���4��s�˲c��}�Ĕ��H>E%��q�Bi���Y����g�o�_^�@w��4�:�Zk��KU��x�=���\�$ �zZ��m��"��+L��DĬt�j��{��e��.]����Ai�Z?�l��n��TG
�`/�&���N�z`���@sS�E�^6D��7%s*z��~�
��A�F����'w�?�g'�ryY�_��G�S��^co1�Mf�oE��� ����i�.oK��b���H�UB��m�J���`�]XX8/pi��w�>�ߨ�bƣ�8p�EZc�r+BQ��؈ܿ�"S��C�kvu������`ǁ�������H�Pi"���#|m@�S H<,��Q���"��0�^������ś�\���<���v����^��l��ɓ�6��QM��">"���/w�.3�og��xJI�I(�ё���iV_��L���T��(�u/�����m�5��X�S���v\��\�|�O4��#;~�S#s b ��/����������\ҪC ��~�8�w#�	��*_>�n/�Ʃ��ݪ��]�^}�+*j�b<�י��i}[I[|�n�uS�4��T�͋Z��w^��B�-������Oz�t���kk��M�����	IBq ���߿�@N���o*�f(>\��d"X��CCl�{�~�G9 �$5���������a-��h��y�`���0⺒�OOO/���nd���������`@'��&�`�(�*Z��߷���<;�{�+�s�l�tЖ�e-�բ"���*nA%Pbj�υ�אH$T�h�]z��� ��(Dc^I{�z��gf�[za��Z��:W�:|�����s��s΅(�ٖ�����'�d�Q(�1�պ��aU9��z��|��!V������ة�DHh�0���f�owH�{��ctl*l���^EF�27"��f�15��,j�T�����FC�ҷi�������Qr	��^�z�B�R�Q�
6M�b��\��M��H��V3}��F�Ȉ��ܞ�=��{�r�A�ny��;��Z��þ�u��slŃXf�ފ�{L�K@ ���)ZT#����U|~ݬ���|��̤�P�w4L&�p��?E`���oE)��WQ�:��l�7iln��B�I�/Vx������u��DUIt|B����KN'޼��4g��Q�!GMZ	�Sj��������/f�K���mx���@K�)�L���Ka�������~��Wc�h�'<�xK�g�ְ=�Y(��0�bY'��$ �5
5�:uoJ���W��f'��ґ�t����aw���o���ob��6'M��,{���nkS�/�&/�٩r�h9c��ԛ�4}i����/+�	��g9�
ǖ�o�sY���������C���^���� @w�q��풏c���r�E�ħ���F�[�б#�ylT�� TJX����}�m��=�� �Ӄa�}�ωKe������APA%��*���r;��dg�}�A�IG�Zx<w��j��wq2���|�n�#�C ��@�v��	3�������}NT[J�(ƅa�hIr�x,�iG<I���&	�g	�1�����5h�9�ڠx�#����/�����{6A��I62R���%�rÙ5�r�+>���i���a>�v�b|��s<٨�[ы�0�����v˃`v���#N=���F����waL 8	M�m��@ �>�����箸�X߾}3+.D�d3�qPn�,F�$=db��<��T��W�O�6�b��cN�+�:��%{\29�u�?��m�|)�C�e3[��C�P�}�]���9�{/3cfb}rd���4lҒ�|�3O�Q����O?� 1�8i��#\�HƄ�n�?�z
�y@��6�Q�p(TW'�,\�������s�����,�gįp��'췞sRSS����A?�ᱜd	�����A�wI%+�`N΀�Ls��Y�Jc/C��u�j���g��g�{|�.�-�Ywf��?�&�H]�c��dP��2�y+���+�|�	2�U����T���-s?�4M��s�F��V��
���W[B{w���zR
Jf���TOG���e����#�v�7΃b���%�(������?�@c�l]�o���UÆ=����V�^�9����J R�t@�e��yEYtDm킞M�D��:W����#�L@�mo�H2���yZ��l��v�	��&JwO�}��> W��aqS�'�c����&��3�3���{	��q󒀚é�b$g�>��=d�*�I����3g��lj�,�8��k}gy0#�n�6�+-�t:S��۱���,���v�F[[]���g��#�~+�ƁA�v��p'�����~�?���|\��vz��D�  ��z[/^!3'o�g�4((��h)qxj*�c fJAj6� U��<.�5?�[;h(���n�q�z�R�qď<1��`v�ubf8��i�+}@�u�G��r����[�<@V{�	�`��#�+�|�����`l�)Zi^��ϛ=�(>ȣ�8Iz�$%���O陮�n�)���#rgE������3Q����� �޶/4x�`}..&�#I�%�>�����6����t1��'u���VR?���l
��Z쟤��ڟXG���׿�f�������ZVv6ε[�-��ė����@q�.gq�.��e�,�:��>P�.�7��sj��QG�8�Z�4 ��S�$ OR���] [�s@�N�!Wp�s�#���O�s�D����X�8���rd���N��Edj5^��ht��[ *F�d8�# �C�sm���;�����{o�!U��!�03�eNK=.��s�׭���#Q��\gKN�[ކ@�����w6�myϝ��M�<�q���g�v�}��<t�G�t��X�L�/��r��`ޫ�=��Ts��C��Y^�9�(L��� b߀�b�7�HP���!�U4Q!G�ä��l�C����wC������K-�X�ed��K��1�+6��X,�6�����{���X�\�24��3:;��ؾ�O@�-$v����KM/��/r�W%ظ��ST�V@��e��1`��"�O8�,�4�� �Cc��ٲ��y_
nm����1G��"��2_��w�s���)[�0��� *a
�`����C�����#=��ծ�:6$�n��%���O�K�%������C�Vh}�׎�]�n+��pn#��%�� �U(����&�95d˜@^��̊
^x�늑�s?����s�'��%�OW$�[�֬�^���3��������V����Ff�����U�v3I}����u��;�9�@�g�Jf� ���Ҽ�X��~Z *u�a�[�S_�6�ޠa-��\f:@L��R��	Yȿ~3(pUh�Pr�+ �HxR�zD��u?UE~3�I�F��"� ,����q��쩨�v�����vo����l�[��0�c��9��쪧c��/���$�*ٓM ����� �{�+,�Ǌt>�������}OYC}���N4��� �]  ����;�����m+@[0�kyev�<Яt��c3��@����s1���"��	��N'D[E/�ˑ��Y��e�}Q{D3i,�&��}�61*"I$��6�OA��Rw�[je�	�(	*"|�ϫ�<K�,��3a���C4��*�~w�|̜l-+EM"���ȏ����:W6���ν0W /)@�@�(����\m��AO`z�{��I1�� b��5Ӆ����Nj�FDD��������rj5�!�d�}c*��Ӿ��T�c�����dWp���� ���MKNƆA��� 6�J'	��%�AS���eGL�=�2{�d��	1�ܼ<���� 젿�EU_�ˌ�(&�}p�+>�K���:��M��u�<�MM��A&�?����ݨ��������,�yK�>�,�b�*�����b�"'��5�ɣ�͡�ݠ�*������Lw��9���"h��;u,%F�e�Gd�C]	M�'�.<t�-]��ί<L?z��鹓Y�vږSis��^-V�TQ�Ũzzxv��+�'��1Ӝ�Z�޶Ɖۻ'��7�_~�f���ꎺ}�t>�`��E��y9Cù7���G�.k��؜?��QKX����E �g�����1������$y����z擩�bg���������#�m�F�g�������O���	�ic�iT�R��Y/����E�E[Ó;�4�إ㑛��Y'Ц���ם�k0��;?{I�����p��]\���|F*�ֈ+��D������6!J��>�V�����OZ�7N\��|n:���>��*�y����d�^�bߤ2� �n�	� C͕�w����������wX�ej��	I�x��m�[���
�`�˩B����AB;�T����.��]SB~�_�&:n���@c놛)0Ԯ�<:u�������9�=�~�	4՝;P9$�n����+�[��_�� �%Hh��I(ğ�����R��X������x�����/Ǽ?��!X�� ��̼'�=�����jK�����y~- �y��N��f�v,�$�l��@���G �c���K�I1xVg��&RkǼ{w7I�LL��uC������j��$�`�����JZ�Pn���ӝ�j��h��qc++f1Ó�l�X��!J�����Z�G��,��rs�J
�2|���uh�KH��e�ǎ	�o���rI<�Ӗ\|4=�</�7����zUq$�&��d�����I�i�/�,�QM�T���4�h������V*�+��^^^�9�­"�5���Z@P�+}j���u",ŀ%��^!g�Q�g�RP�B�8ZZW7ő����Ǉ�� 3`��1X-n@Rs��qVGi�����9h�7
�C �''u����z����(Ҙ��`���X&P"�Nr涺v� J!Űӌ���q�-��sj0T������Ek�D� i_s���2�ŧtj:*d�G�6T~b��Q���?gՒI��V#.�������L��8�*M�e���~�B9�2m��W ajYKɭCm�E=��!�\|}��8
%V���(%9Y����X\����)��V��7�HȦ]��ff��x���eC���;P@��|\\���#� ���$>�[�/~���=}g�P��h�}P�t�˱T���Gۂ:�
ia1�S�0�(	��g��1f�P޳`$�+��U�Ҥ	`Q�B��V�@Cb
���ݍ�����eE}|3���a �NN7�=�$�>��	G�ړ��|�2�+P��6��җK��2��C[�?^�)$I���p��X�,�q��E�J��`�"lC�#��K�Q�����s��r�B9�[�<}Q��cr)��[���L(�^X���e���������`�x�98`�~�F���&9j��������+�U8M�Jk���M�O�k������K\q	��"RN�7�q����ry��>�(g�1�<l,EE���@ .�X3�'r�.˳$O
h��m�I����z�8HBq8�e�yqv�J�̓��8��y���F3��x���'f�誐�l������M¶���E���.���깜$���ԘH�?X�w+�x8K�\)\�5�f��R��º�z�e�`$�J���`]	T��UH~�����mh�Y�C�"8vK�͛7/����{��Z��Ƒ(5馔�3h_)~�AJ�Ԟ��W6�o\5=_���<'���z�_e�
�>
 ш�v���e ]�%I=�J�ԙ*�� ��QK��`���L�)c��}���#0�gϞ���}hw��E��e�z4�>lVPT�T����<���d��}���5j��'u���
Hx���B !fJm��=���/YQ�Rm�%�6 t:&&�58�apԏ��:,T�U3��r�1}���>G�w��,��m&Ů�ӒQX���뿱Ġ`w���N�����F.�9��jD�� u�3�;�&Q#!@��T���tM)�$7��Tz�zTh9݉�(���>�J��ț���IA����:���P��n�>#X;��Ȉ�_��;�i�i^n��cCA�u��"�1��~�����xM%3<:������C%�c4o���9�K!�,g��+�`���&�:[P�^���||��$4B8$P�:��c!8bξx�}���y�H��<�� +D�yx(d�@�٫Zda4���P�$�r'J�_���.�qT��'���/�	�KN����$�٫r���V��)�Z������ؤH��,Z$$#r���n�%���rw�V��DZ����D�Ĵ�l�L��bB����g����|��s>���<������w��s��~��v)UA���X�#���fQ_E��C��n &��m窘'����g�yJu
�:2��sT��8���9έ2Lb;����̝�~�>�gTK����XB(^��N��WC������I��y�7��������w�^hXx}P��O��O�J�R�Tfn����/.�9r�MR<��q����ۜ*��8������:�x9���!
⍿�_'vumhA�N�������:?�~|_C�!�pg��j)5uL\X�I���\X��U4��b�cc�-�� ��9�R���FR����?���O�L�� ����M����ӻ��,{=8�2�L�AJC7wE�B:rhY;�Z�~Ȅ�*��m؎��t ��-��DW���R��C�Σ�?�>����'Ƞ��h�{���F@Bݗ�2a�����6'~�ę@81::
>������C� �`X1n�����f1Ƹк����t�]�kH��{����U�[�������{Q�4q��4�
��`�Ğ�08#j$'|A%+	������<o���/�� |��� 4�����^Q��p�Dۛ���D��'{5��۳Q4g�6}Лm�}�S����/=�#��։��,*����?�8�*pFH|]j����/�1�A�{�2�0�$�-B��r�L�#�+N<x����t�%��|���N���tJ�Jc�n�ɚ}��f�NDg�,�R_���A싿`�_a}Y^�r��S�F^bwb����/�C}��%�{!?{z�= #	u��Ŭ�䏻N�ћ�8���ȗ�y��sו�{I�VBv/�.˘U������_?�h�}!�����?u��Ԗ(/m!�}��ұ��N�o�NO�^����؍�Y-�YK킓n���DE����t�����?W�X����Oߘ=z��m�I�p��I@�N����m���b��0N�ݔ�R����Қ�eͰ�i�C\n��Gs��L����ٱ��)�����N�����?��@���p�� ��t2�v�9;δ�|M�YOIh�,�e�S���vDV�_}M���1V��|�Bu���;�q��kS��ZsZv�'x�ui� ��T��m��� �U�������M���`��'o�s�Բ�Z�c~
�qw7-C�1p��;ځU��wʁ�am�{,�Za>�wxm�}�S�T�ۭK�y���Z�%��5gv=,��11ۼ��cEi�3-&Bы���6�¶paa�,����Ͻ���,N����&���@���$GK�єX^Ĕ0PvL�e_�k��<��C�x �^�J�<&��I��ݗ�x�g���0��i�=u�W?z��G/G�t��:Ůd/BW�v<�g�f_�5 ��:�(wʗVO1��M��-��[���q*Ԛ�(J��H�0oE2�k9��hn�DW�.�g��u���Q���6��2ls�]`X�[׀t8}Oؤ�z�Ʀ|n�`G�Lwp#V�N��E��Ս-=>)��W� �d�0�.X� �a� �v�Ttk8jI�&)�a��WH��ݰ�n)����Vm1�����g��{ya�sn�@N⩧�����K�- ����͍��?"���y_Z�@O�NM%>y;�zVP�;�[��l�A�V*�u@K�]�\��<�̞�P#� 侪���2
�V��勪�ϕ��P��Q�����'~l-5���o��!��5$+ ����y��V�5])�a�3$8���^�/���P>�#B��w����h��ZW�LI=\#�nO�㈛ۚӓ�d��ٛd��7/7��oQ*1�{ -������\���ȩ��?���_��K���cuC��Vr��^�D�Bcu;�qq�)��G���� ����Er;����� z9�R����J���WՒB;+".~[S�|Iuss��:��b�C��S�F*��N	��5����ֱ��؛xf��c�`!,uu������A�EQ�	�<
e�i�L�jCtce$ѭXe>�-- R�������-�N �2l{U�Hy9N[\\,!��'��Ù��`0�����W��gX�Y�S�1A�usí�A�m��p(L����?��gef֟���V+v����j}t �.D�ܜo�8���e�Q�r%�~C/;.�JZ��9�>�nU��1�cQ�1���F:��A���J�UŐ��������9eG�v�Q�� ���2��g����v�j�--�7�q�JpI�
���
׭���)�i~����6����$���p��Ļq�0%V���%�g�����#�P8Yfܱ�@d��cͤ������355��~̖�J�<�H�5���7C����G��WX6xvWUta)D�����wH&UBo��m
��\0h��]x@D�F�_��5@�"#-s=���yDN�at8�뷔��!8 �cqa(�EF]�5Pj�3���(JMb�k���3��[�P�KSqP��/�J�쵥�|*�ߤm���1�%����::��}�e�	�!���ȯ1��m���T�Ǥ�\o�b��"l�<<??_1����PC�a^D����Ӫ�+�rz�������ZW����(#kE��ܯ�g���,m�(�=���������%z$R��E�͌,�/���/PK   '6X��g)�
  �
  /   images/c1fb8ae3-abb7-4800-a199-c8a1e0562abd.png�
!��PNG

   IHDR   d   B   �s   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  
kIDATx��\�k���߻��d�dK�jA4F�H\BK��N?p[���/�C�P(n�R�?Ч�ҧ��o�@����UR�QS0�cl�.�lY�W���jwgz~�=������������;s�~��9�s�LBD�O�<�D�B�0#�R)�L&E�\��j�*����$bϞ=b�޽?��o�YLNNv���#dvvV,..�l6{ƶ���,�;*��!L
�{t|�ɓ'o���v���#d߾}��ݻ �;��n��������W�92H��I�z��h7"G�Ç�����HR^V�h���e?Iȫt~���Gt�#�l� �aQ�>�����C��m6�����F?�jK�Eİ�~�O�^����/؏���m��\.W&���������!���bbb�P>�o�V�#D���������
gΜ333�T*}�:��'��h�u��3���=I���b��	D��X,b���v!�o�p��
>pR���={&8Б�G�8u����ܿ��D��d)�N���3�������;�������"GM[1�] ��1��$ #.;�|�����z����N�:ձ�G��+W�xvg�1�T�P�����uk꣏���?�޸q�#m�!Q�sB��	�2D�uP�7a����;�B���MY��۷E�!�<��!��aw^y�uw��!��:>�!�t���'�����ѥ�·��"�Dx��dv����y�cc��4.=�����vD�t(��[YY���L:$ ����d��w���&����(��P[4g~��='d���.ҹW��&�v >YU�&�رc"N����0��r�:�P��ᡡ��r�cI"J�&vtx=ச���?9��[u��r�DMOOSL� cy �H�S͝0
�F����ˁ�V'����>H�#�0Hm�I$(��. �	��ras j��J�!���_��x0�u%5�OJ�*"0!���h���������d�C'.-/c��*O�m�ȧN�C$�.��:�UҖlo���˷b��ϋ�J�a�	�H�(��!��m^�0����͂���P�\I��!0!��8#T��`��ُ�2�F@����יt��,����BH�������>̕4��k�@�jnb����ٞ�(��5���`�7
�)!L4�
��2�'�G���SL 0!<;	�Ӹ�L�I���	�t�2Sf�~eɝ�a��`uez󃖄@l��4��4! :�7��,��U�&�B����4��.B�d�I�m����u����*�ج�;o��@�����J��.�v@�=��>h��@+�v�����κ�iG�:.!~e��< ��?M�t��ۅB[��݃��&o��|>��:jbB]uBM����9��J��!rX�"š��;�{����G��6U144$����V1�׮]���T�g	Q��TWu���ctl__�$!��q�������c/^������!6�����t��9}	�"��t��gGVΓ�;$%����~R}������{cjjꗃ��� �7M�����oY��3�.�:nCԭ��N�w��Mˉ������$=��e�))�f�I��`��X�G��g"�W�.]�300�aGgY~����_Y��� ǹ��s���]�X^��xNrT�K��xK�V�U���1~�lB�y~�h��Ż���;`�k\7�Ћ�Pw���z;�M���8-T�JKH3R��dB�`9-Bt��mZiK�XH���u��#=he����K~�/�-�D�W./���4�W$;>�m�����x�r@R5�|n���!����!��U����9�V�??�mC�H��u��W��Z�F˄�$��i���v��V;�����*�<���cx��6&��sq���"F�P��':�`?��OB�#BxB 8��<[Ӳ!��� OL�#�-�	���dI�+�I��ȟ��6ꬲ�V+��2	Yu�/Gk���5�!�kE�C�:�WiYe�yΕ6��D6��m�0G����=�>��C(���5ǳ�Q	Q��F]U���!->Hû�ePG㍫?Y��5;��S	e��T櫵r��)�#B��$�S�����E+���)���-is��CTP�Z��~�����6|ޟI�*"	��B_��7)��ׯN�<�/����9�8j�!�mB�0��Fj�-L�Q��8z�lI!vw�w�f`qH����fg��ŭr�r�5 �~��Y1���������+u \k����u�a2!��N�:�\�{�m�N)�D<�X®�˗/�x���m%>�QZ*�ga"{�&�JHPpI

+�Lf�}�K����و ]!!rX�$���Q3ݽ���9����SHR�I��%�7Kk��d�jB�3!�&��u��&�p�~�\i��E;�ʌL��l�I������#5C��l�oT
��m\;�]�����׌j1M��BB,� �
��8n��{���!�n&��Hㄔ�ٯݲ7^v�Tn�qJJf��,�?	��{6M�]��u3NȾ�����<!j5���%���p�-�M��m�	+�z�R�,��	I���<dD ĉ���P�\+���:�nW���t	1�.�T�R9�n�B}	q���|������۵bص*�
���7K�X=v}��P	�?l��v�l��k0xO�n�����Wㆰ�v    IEND�B`�PK   '6X$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   '6XP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   '6X�.m�Q  �     jsons/user_defined.jsonŘ]o�6�����3~��H�"@�I�]AARd"@�\�jP��l�i#Ѧ� ӅaS�������m��\�Ⱥ�k?Η�+�y�յ벩�����ug�G�����O?��}�w�]Y7�O��A�7�i�����m�ԛ��*�f7��@��8����ge��aRF!�1�h�������y�nm�r��M��Ci�oOq!!+ �BZ $+�qg)fV�|U߆~���	z�����.��	7Ve}V�&[|�����\�*����\U��#���ö�:�v���/]�Q}V\m�2���Y���ߗUhA��9���r���]ӆ.�b�vak*m\�ԧ�OWoN���4��t;l�����͟Q,cY�ҭ�&�%c,O�\G�tLITg�1S&1ߞ�_C����$�uh�A����Ke�13���L���pZ�/q:N��%�Cǒ�i���q�XP8-��,�I)8�� ���]�:�(��=]Ʊ�Bi���ƲB8��O�h,,DҰ�hOp���h*6.<Q�X*6.Z<Q�x*6�_�D��X�N�,�H�q�Xc۬�Bq�Xc%Ry�:�ض�P�YO�-�H�'D<Q�h"5./<Q�X"5�.2Q�x"5..2Q�D"5h�f{����e돡W8��ؖN%��JF%�C�	gw㱆� ��U۬\�)�0���n���������궎"��>���6���y��O��Տ�^�\��r?�Z����w{��'6��;��k�1�i�x����Х�]��~�S(�⽾u���v�
_��V�;�}���+N�t]�jv�ј�Ʈg.�>4��F�jm<Pk�<��Yf��x㙷Ф�+�}��\�5��@Qc��Ġ0� �>��=6J� E��¹�P���T�X��x��9�������_E�x��\�\J��9���ZWGX,�PΡ��_ �%#��q�b�8'2u�mh���P�s�C�/@H�q~q���H�nۦ��XR�%?���� VK,��EHr
 �7���3g
�����WPs;�Ѕ$�/�ͪ��ն��a�(,�@��%���0�"�Oն�^�� �e�m;���[c#(A����T�I����(�*����BH�� 4\���>9F����.F�)V�����	��@%�@#�B���A��)^/������ػ�G]V���a�,�o�r �T�X�(�����Ea����)���"�5�CBE��{%��J&b�y��SH��{G!Sl�;g�'����G�8�8:�f`� �2����MO��=���r�byvV]�'��U|��in��i����a��!�Z���{��PK
   '6X137=�	  2\                   cirkitFile.jsonPK
   '6X��(��8  �8  /             �	  images/02932828-f6d4-4923-89fb-67d65ebd103a.pngPK
   '6XR�\"# � /             C  images/16f29068-8fa2-43fd-94bb-aa3b1aab738c.pngPK
   '6X��g� 
  �	  /             �f images/4f5a6b59-a216-44d1-a198-112719b334c8.pngPK
   '6X�� �f  y�  /             �p images/96fabd4d-0b16-452b-94e2-688cfcbce531.pngPK
   '6X���5�  1�  /             �� images/a437e5bb-8d3f-4b3f-8093-72e2f97ca498.pngPK
   '6X��g)�
  �
  /             �l images/c1fb8ae3-abb7-4800-a199-c8a1e0562abd.pngPK
   '6X$7h�!  �!  /             �w images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK
   '6XP��/�  ǽ  /             9� images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK
   '6X�.m�Q  �               �L jsons/user_defined.jsonPK    
 
 j  R   